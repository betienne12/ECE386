XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G��܄,S�1��W�0��S���w���x��BnF���/�y����)�%@�{�����B���7�ӥy�r��cא������q>|����Z>�/'�_eOe�*���
Vy��\�o�.|}�x{5�]��\:�L��)�>k�b@i�')/m8��e����ԭ6�+-X"�iG��FN1���W��ID��I�B��[��Wa���Pl0�~�Kh�w� sL���2��v�F�v�OE>��Y�3������32<��wkD�D&H2Ŷ@��]s���r�`iQ�Eū�vx���/���&�Ԉ�iܰ҈��fW��崵��9�T��6SP%6L�����3��B�fcB]��K��)l��9�Tw� 'j�@�Z�1t���}�`(G�%ގ7�{��i�����^cL*��#���[��/���_�@��&tܕ��gﶤe��L�Y�%�>�]/�Kt�{XSF���{�3����V�f�u�X��ѐA�,��]p<n�.��@@4l���o�x-�O��R>ރqԠ�,Zmy�j��d��5&�9�s�/)�-XB��4�$���F�N�H7mS��ޢP�[�D��a�@�W)��mb�,S�d��9��@z�F vs���/������E ��3F�5_��}:ʭ��t.�Q���6;#&��ռ�	��Ӗ�"-��SM�����T9�OBM��&�����#�VWk]�P��um	�mtPd���
�{��0(I���,*:�/��#�XlxVHYEB    fa00    1ca0��
��;x �Le�_��1!룺ȌѺ�iV�}��c��25;��B61@:9_d{��چ�LNu�x?Ab��,����{[:�!����+g�����U�a��?k6OƵk�Ҷ��G$RF���q���M������ԥb9Y\�R&O��m���L����_gؑz�X�7��أ���؅��-��#	��{�`&Q�E/!��h�D�)f�	�~6�T;��C�Y��Ҩ��5���]N2hN-U]��??G��H�:���)��!�}�$ɩ��K��8��t��GWI�&���__��괈�-n�@��� Ј5eRa֯dq;>h犙ِE?��T�T�Ҥ���2��']��d�u��#�~��c�e%������[_�x�}&���W�W�Nx>�,�kA��&D��עF�$��Y���|���nǋ���k�>�+\���&�ۂ���>���r���Ё$�n�(��S �����k�_dS�O�8g���$��aKT�ؔZ;�_������T�4.ƣA��Ց:�|��hOߑ;�������E��Y�ë��}�&����͠ӆ �sF���ʄJ4����{1�;���3���M��2P��Oy�4�b� ��G�`�����ƁiǣeA(�.�:4�$�~b�H�G^�~*�;7��*T�fˍ�ۇhY��8�D>��" �dQ������xu� b��}ٰ�����X�3��Nț�O!2u@�i�^ ��5=��KX졄����y��p�?���>I��C�� �{E>����A�������d\o�E�%ȏ//T�X���VS)��L�A^/ش7�z����dSJ���o:P�@���A�-|!C�(ѣ�4���O((��x�X~�U�R������^=��M�]F;'����O��������n���>@
<g���zY8T0y/wT��?/1+�p9���B�.����#����ne���C�"2.s�^�����enooc�ү���!�jJ�u���G(>���X��G�'�K	��zM��W���ʨ6Ku�d�C烬�̜j�á���}Pl !4���`�[@��{=	�?�6::�%b�Ƽ_�HU�DF�V%���Ƨ��:�?�6����1Yh�ܣģ2���޳��7�,��� �M.)�	��L����{$��O�.ZIZ��Hg�>�U��l�s��U�N+��7��KǺ�ɬ�> !dP
��2�{�K��HG����~��G>���6z�T�K��[�V�\�l�+��Y���)� ��o2�}D������#�Z�|�R܁É)� ��>�e=!���J�6����f���ֈHWf��^�Qnւ��+�4EֱK���h��
�G���i��:�8�$9o{;�=/_�z�{���hg���7�#�o\�Ʉ��e��2�U�'�J���k�ecV�+����᧕�^�zIi�am:�u��Kzc	�V
���DC͝V������v��x%���3���Q�<_4.L>U�#M0�D����/`� �B��#t�4��~G��|{�h�>��l!u���B �F�엌�@!/OµïT�q�L��*�ys|�F��]�����)�vܤ|)T�y1��Pf>.��i���$L�(D����6��:��5#�
��}�-��B��W�hj��.m�ވ\i�]���Ž�d̸�4(��±l�����=OQ_)	ym �cE������V�{m<@�������	rp݀d��-��u�NN�	�N0��ߏF^��?;���ߠ!(���E+E�Ed������`㴛]1Y�֍Vq5~������:�-�oH��b�[C̓�*���L��Q8��Ӭ��z~�*677���q�k�p[��͏H�J�J]��O�N4-�P#m��`Æ��=����l�!b�4���AIY�t�:�����}�4Px�9W`O�]����Er�~�	n`�N�OqkO|D��ԏy<(�S0jD��x�c�z��J��o��q�Hӑ��{@-�V}��#�������]b>���^��2l�'� �&N�rX�5hq�)��D��hX}��+Dr�Ʃ�o�l�I�;AfI96#�\�q�����C5o$��3�T��Ud#p���b'1���K
�~	IU���7ό���I+?������X��H��x+�'�O�S�G��/I�~�X��K�d�>߼O�ܨX��\6��9Q�l<�gi����=���&�/��ٽIE'��<Y�̥$�J�9W
�v�''����E���g�	^Z�զx�(rO��ّ���9�i��H��gQnH#qo�ɕ٥h��93Ꚛ���*!R}�k'��9�=|��W얠�8&�O��)�q���6�o��\�8�~gR����l?�>�1C��� �.3(�o�1�Gn�n.��*�����"�͚�Ι�������e�� �f-|�+�nE��\/1;]6{��}�4�۩���*뙕�Fx��#l�HI�<��$�,^+��5n�fJ�R
9��a$� Z�˙OR�c�B
�Δ��hMy�CԹл���Z�K����յ��/�l�b�i4F�O��]?Y���έ�Fܹ��`��c&��_D/$&%?v�46q��X��g�s��59�|�3Ո�K��&b�z ע��4�́�#�н���	�=��j *�YU�b�\�L�;������vC4a6�Y6�d���ej>�
�c}^!ڀ����t�U����2sm	@Q#�G���7�m�+�H��m����x�`�_�,"�x��N�|��Cffi�������!M;|OpD���/��NN�.[b���-��rP�k�^�7���w�D]'����^��ǈC|T��Ⱍ��Y�~�wC�t�mzw<�o[�O� ��4�7�(2������>^WK�de��x+��{.��@�g0g�:%�c�cڮ#��N�af;e�ɊJ�a�C>T����`�
յ'��Po�K���6)��E`V�u���P��2ֆ��_���sڌ�F�ݙ�0�61��	ob���ΰ_G�γyL�8��7��P���M�(E�/���<�ő�>�sg�F�ܜ[̶s��}�,�҆�J?6P(oȒ��!o�8�/˭���O2����yqy�������L�XZlFϨ̉�����l��n+���xPg�����g��`�}f�߬�{�r0�C�h�Ғw�&����tX��<R[EÙ�8%��&�J	���3�w|�J��ًA`	�F����z��^q g!y��z#Y�^����4"�^�"���l�RJ���@�ÙjM��`SX8��ם��#��sgm�j��~ɾo��+�8�}_���ȉ����W�$����2�3�((x'w���L�n*��%�a��\[ٕ�ި�Z� ��J�I��[��4���S��6�vX��m"����d�R�67p�e�����O�N�E�?E����=g�sP+�%e��2}��>hn����Uc��#�G�	-c�iuL2|�<M�����n�q̭�c�
}�jt�:x�����%A�L��0M�)��uQ?��,9z���2���M.Sn���� ��r�8�l �.�`�����|�Z��ro+��Jbw{=�%u4�����5���H�}�k�~�R${�(1�c�ƍG{v׊��﨧�C[�4ލ;���B}Q����ՠ���X�ȶR�f���ŷ��C#>W{�}��dш�қeGLjyj���{.$���S.�?���T�_�<Z�*��;� �[�,�
3ꨕ�����女�O��.�X"�M��v�ȐiCS�*�Ո��U��A�Г_���>Bͳ`�BS�)KԼ�W��@W��sR�Nr�n��8f�rۜ`y!)f���k"=�Na�����_�`H���q��u�{��NU����-y�B��;�4�c9���H�A��#Ο�ϻ�Je~����v�cg���v���B90���KihS7�5�y���\ы@ȫp�D�GE����Ō��dD�~�������Ը)��al1��3�-�d7 h�K��t3�u�}���1E��49��7ݩc�����.>\DUD /%�π$����HD�[]�~�z��x�9��a��!2��u�ү�vP�`XU��vh�EK�<A}/�݉��q:+;t�:�9�7kܚ���R��k�ːOb?��%\_�:�Qp��a� �����h�d���]��&�,���l�q!T7iү��6�g�%F��{|Ż�nqZ�4��5���/����l�G���۰00�{��-�"��r�O`Z��Y�p�v[Y�3(���"z^9��t��\�5����{ly�T��W����!<�jtȌ��=(��i������$T6�g���ΎF&&�`���+�}��#��
�*UR�B�����C%.�
���r؄�Sxt����SD
�lx��=n��!z=|o�3q��A��g�#qہ21>_���y��&��.!�g�����(4��sʿ]�Z�==ʋ��
�����J����|4x,�^D>���}v5^ �-�s����Zn"�C������u>����R+�*��&����D�n��#s��ZU���D�ݿjj����2׭�; �o�y~�rX7 ~�رY�q%��D����t�
��2��P�� �<�C���X�[�e���kU��ۮ�M�<<I.�\�cB�c#�&~��.e
��]	��)k�uj������{p�-�������ȧ8�0�v;�@�*�lkf�,�
d�|�!��&Z	����n�> ��gz��È\��\R��=Z�-���y�\;uS�Q�|�OqVh�E1�UT�vB:��7:��[�sõ�,�M�͜��:e 6��^
 m�~L�wa����,L�}�Ϊ~q��&��T�+�=N�K�ރ�u�T=I��v��F�B�=mP[i*�>�34�����������܍��ZX�P�
:t�Kl)Ɯz��&�PK�o& ~��G�޽]��`U�i�\Y���� �ٺ*z:����vp� ����>� �,�+���}�����'��F���n*�8�f*���`
M������3G>*2i���lǪ��ڛm�)�d�Q&/0e�Cq��TS؁͞�A��`]�v�]BNn�Z�����hG�eP���M�_
��{�XĔ	x����J?.hދ����r��mXFx}#�:Fm"��0�6��Z+)�i�����;�Le�8�LR�be��v}}�������F/� h������q6��_A;�W1ޞB���l��V��Q��e�� �H��yv�`���e����������T��D39���="w����gȑ�@�9����sVu�r��1|����[��"���}b&��� q�A~aZ2WW�H�S���Ų�t��>�3�w<��C������G�8A�V��!��M��/\����#���iP��Vc ��b8����M,0-A�6C~��?�-<�d�FIIea�Ӽ����𒉴�� �����a��aB�m��N��� ۮf����ِOqe��g�U	������,`��Rʰ��t�Xjܮ�2H���E���W/4�>3^��3�2���ro_FZǒ
'�eԔ�K� [���QR�?��ok��������M`I��i��c�R��'�F��}>_U��&�'����If�Xpw6�E,&	=��ހ�Ўa"Ȗ^
��iE�1!���I� �`/�V��<�!�h�Ǎ��e&����ٓ-��"���2���%�����gN��va#ףK�}1��oL���S�O4�>S��<�F�e���ٿ�c��o��`WlJ#�m�)���-qHd%��ڱ������x����j�g�'Jxx�%�̋[R=���j$v}$�s2α�H��>n�����9s�b\I��d��P��ՁuQ�/����aݤ�"�U��)I�ՔAm�H����d��7"S��s �?�`���ly����Whq�lֺz\���f[-��&��g�N^����R��-�@�Ju;Z�	F�n�K�Q�G�OJ̯�W�m�@�+/ m����V!J��h�ċ���)}B�P��JT�-�;M����M��wG�G��ݐ���� 1���!e����yGΥ\�G��(Bl|X���`R�Ƃ�G���]�K^#�w���xj�<\¡cf������)�Sƹs\E�ܾ�e.��{s��;�_N|$�&Q�1y'3)<g�vi��E��a\�D��q�$$�	n��	���X�l�"��y�!�Û���R �&�U�0d�*z�oa�45�G���}��q6�MO�&�S�G��_��'5iP�(#��D�X9r�M9ެD̀n?�]w�^AxC��+����N�ZyP r���r��1U���"��p*���(a趙b�,jY&��_��QI�AI5�\�2��@؃D���B`��]����o{k�%�d:>�QFfJ5����&��e�{�!�$]a\l�7����`��3�K3z$�ǉ�A�6��a��F�����
u@a��#U��*��:��t�߅z_/����x�Dy�_�R�rC͖�֫�{v}2���}:'���a$NG��YD{,�����2�Dqp�Œ0ՖS�����5
E��~
u`ۚ�,�f)��2��_���Vf��l/���nx71�����
=tah�����H����,��G�7�V����~����R���)M{#�[Iv;K�r&+���h��FAm�Z����>2fK+�:��r����w#/�F�х��}Q���x�e��\_��/CU{m2�}\����˫b�=�_����:D�
����^F���
(���~�U����7�08��u�f_��A7o�!��t��	�n��d��64�o�_����$��
d�(m�ͣC��ok{X,Z.�j9��+�Y.P
��Y:��_����d>H����b�XC�)}m���+�r/�tXn���]QypC�tt����
Y�V��zǣ��D�`^�%ҐTF���.	���`�329�ױx>�������.��a���9��eE�����s!V�{zkO��S�e�؇Ȉ`fѠ�tT
�wW����CiR�-6��4N�d�ذ@GfVA5	�H�݁9G�Q�neX�w��N��?��2�&�C�¦�D�%o,~"�?�l��Z�����^&@������	�ix�\�{N�\inb1-�XlxVHYEB    fa00     cf0X�0x꼅:[g	n�
;e	L��4���
�����ΓxN�
I��l�R4680�s-����+8��ڳ�4
�}o�w]��'�u�"����TȚ�n�W�U�(�˝)�Z_�2�q�����d7[���w�^/m�	�ۅ�6�[�����:�4�&��Jj� �웂�>N'�#��P;�G^\�pݕc�'Fr ��#��cCX\�p[�B� bz+��kqp$\��)!lMZF�� ����k�-����'y��yM��u9���*kwˑ���o��V�a���x�gK��DY"��HP�hؖ��K���(�a�C����D}��ٛ��!��6����ݶ/��Q��CUl�8���2�25ό	ލ�(\i�UNU��ǫ���qB �r���i3�J!S	Iy��M���T��7D��]v0m��U���b����t$u��!7���c$����:�nj ��{�gv\Ѻ~�&����;Wm#
}i��rqg
���̏�����wFr����vB,�\�����&(̹�#w��FA�6?�Ι�ߙ���$�%K��Y�O
?'ʋ~-i;�c	g���B�^͜�11�ȸ~�)��x��qnz����/k���p&u*�	�C��@��t��d�	2�R!�����*5_���%&�%�*Qi��o�_�J�n<��S=W�����h^ڲp��Iy����{�FRAt�Tkܬ
��������*gL�ܤxuQ��h3Q>�2bR_r���N �
Q��b�s~e\Z��A�:����R�x���ۙ��"����b��4t�A.9|�sZ�R��P x�
 ��Ϝ5 ۊhԑ��o�q�0ޜ���Р���^p���xʰ84�s�1̷w1�W�ݥȳh�񭠋f"#t�<�т���s�,�L6FC�mO��u%�3�l���s�i��D:@pI��ϻ9���х�2g̠A�4|i�T�H�N
���̓�!�Cd�~�6�:ORy��T�9���V8����l��R�͊�	u_��_�c�Z�c;�J���� ��UT�b���G5�o�?Ԟ����*�풞�c%��N�qq9�@TN�`{�`P���c����\j�{g���VO�q|o�Q��"��A1i,�@N~s�eFX�_�Hks�`6��}X��N֮L�����W��n�0p�&n搎oA�/ä��v~�́��#��;�i�X@C��pL����I��i�#�F�Z�$�SF󓰛϶x���E�-�y��o�YZ��C�j��K�ƕ�HSJ�Ec�@�����ed��D��}���lK�Ą �q�T�C#���j��4k��ib����_��v&���EKt����c�t@����L�����f�9W+it���A��´(����u+��>�dl�(��ه��O��1�$��_���4x�VF�N��y��X+�8�%T��R�F$�ָ-��E̓��~B�ɴn�9+�7����xϪ�;����1��eM��𻬟����	�TR�}`?���R㺝���~���~{]�b�ƥ�[�&��k ؿT�^��}�e�������<!�L��9/ZU�BN슩e>��%zǘx�o`�L��$��щvr����S�*O��z�Q7�VF�����׹޿o j����.�Y���cn{��N	@� ��:��YI�n+��7ם��}�Q?R))�܎�l&u����u_9��ioS9�\Z�:pH���N �C~��(y�7-�7� o:�J���&�������B���/�)R���ZN��ڤ[t��Y�r�b�cռ��1�r
	(iyI¬�B֠�d��V����5s��<OE�,B�K�\&�,h�13
��>r�UO��Hs����"\,:�f���ŇU^��y����b�B�HDՆ��B۩���˴5�\��]��0�Z�������Mn�Y�G�!�7�'�~Ge��y�A�IC�v�g%{��q��4we��p��R�@Z��eJpa����������]���jyם� �7�Y���*�sq����i7S]����{bQ&�p�%��mF~����"��Ќ��"I'��ӀMe���F(ͧ�V-���ř��`
[.�����U-K�G@.+�d���/���7���M�,>%�k�xd�)�IX&�y�7>�͑�Q(\"�Oy"7���(�b��<v���,&S�P�b㷭eݶe1ToR?��+k�p[Y����޼a��6TP�?�[	���`�l�b�&���hV0b�Q��u�"��}FY��*'"�f`�n�f���Yh�3�w����� ���Y���&(f� �f��M8�J���+v�N��\`1�S�����혟��5��"�E�~��׈�*/��$�p�6I�Do��?�������B9Ձ�&����$��z-��������Z�苭�ڝ���N?��u���0�m�����{�W9k8I"ϛ��u}�Z
�f��$�v¸�I�����UAA(�y��&vϠ��|/����* �p��I�-�"�D6��h�Z�6��Ǘ+��#��/���k�[\���4���ݬ�?�v���5�:ʉ�7h.��R���Qܑ>�1�jG/t!�H��7���	�jd�`���D�.EJ���m]1��ox+2�6i�}����.�RÎ�92#��[�w�4ۘ���u�/�.�:�c�Pj���ȺNa�ӛn�k���.�am��%Y��π�b�Ȳ�=�+
߹�N�#8zcJ���\9QԳ�-x"�Z��(�?�I�tb
z�s�]lå��y�⯜��Z��C�|�����W�*��>����i:vt�c�;\���Tִ"j��ނ��2���8U�k9�l�m�;S�O1"���u�xc� Ǿ3b�:��ހ�GN�Y�I���`�-�?����}�y�<&���I`hf�R�<i��É��������:��u�ٶn
2p*�s@���D����Bn�t[��JI�լ��T{����W��_E�z�����7�+�YD<X�5M��h(*�χ��!�A����N,Q����KZB�	H�˰�+a o�Ĝ�	s��DkCU�~�q�!��Nȟ�Z.��3q����:`s�X���yr�x�<���d4�+��lC�)k3@�7�~��L�*�
(!	y�7��\��R=�3!�����b���!�Tn��~)��"��
��V�b�I��D<Իװ��)Gt�U����wX �_��Qae~���(8��	E�q�wA��� XlxVHYEB    3981     4d0�!��d0<����Y!�5�−jtAދԳy.èڷC�;���:LpDb�>����FT́��cQ�GT���hnҴe`������7}'���qtԲD�۰�ͻ���3F��Ql+g�mڶ+�d����I��4�(���q=6�J��"����=oW^L3�R��)�t�
?@�y�Z��N�'ӕ	41���V�?��;#{#�-f��˷��`ޙ@��?h�k��q�XDuӘ���m��P5�1����O[�e�ur�~hu�߷r�G��}��0�g/P��:�ȧ�?xAWF�ҹ��z֋�a��ޯ7TN��t	���L ?@�t�\Ì,�Ja�����a5cm�"��E��q���j�� 9�l� �l��c��W����qo��V�Å�
G�I�g�b,:�p.��>����ʘt�����	L͒YJ��ݾG[��/���g%�M��Ȧ�	+�
To��=v��A�y���UϷ#�?�8$��x�+Z��d�|���e�}�#�_0�:����FbX>�	Lm�3�����w�V���@sJ����J�L�E�Nq�W0RW�m�Z�~R;-�4��y��;�b5\�3�
�/c�����:>b%�;�e�&��(U�O��&.Y��S߿�.��zu�d�����C5eiFqel8�-��^eR�\��H����.�E��7�^G�n�0�� xTE�Dl>����n�O�������� s�� ;����n��dٿ-be!���tuC@9�Ǳ<4�}�}��s�խ<*ٳ��bD�e܇+R��5Z՛�w�fo /�'�&��h�N�Tb:@!
g��Hx����(c�sJ�4�_��e��NÑWY�1�y�O��8T}7��=�&�Ju؝5S6�h��b>ʷ��Z2M��k;���GE�_�O�	�$[+����_�ݻ�����=�����]�e��A���ڟvJJ2ġG�x����F���G����N����}�Q�>��Mo<���jl�{��~E�m��u�Q�O���'��L����)՞#�v;��x>����'m�Y��>�AO�+��"D�o&�2��t_���|��s~��� ��,���j1 
k�f��������ݠǘ��΄3�GTa̺݇8קA��,�8x�vh;�J|�o��L�p�8{&d���a]j�I�z�2KD%��ss~1�^A6�!U4߳�� P� '��Ō�.���}=ii�,