XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bh�T]᫔��p˄���W���.���n������9%�����*:��Z����i�a������iq��v�P�ǁ8��\�J�-���	X4�Qz��&���a�Oߺ}��[����ƃ_����M�����Ls��_xK�p�r4]��{��O}�����x�b�`�㾶[(N��%��M�EB���v`�>�6����9o:h��M�~=K�Kevh��vҨ�JGF?A<2	!�l.�{�4"p�f�3�C6��d�5����V��@δ�<��	j��oK���?׻�y�[��}�Pnx������lx�	p�G3��$07���
hV�zO�7u!�n��f~&���t�Ah�g��2�e|�q�I.��s��#�v������
Q�J5�k�Rǐ�.UA�s}\��e�B	�|mq��w�a�� ӻL�e��6^�q)��N+掜�ʃS����ӆ�/�C������*�٤śn��0���&{L{h������jh!���c�5�M"����?�)�/efa��B�7�e��A�f
*��@�#u��(ӗ����� 	;�:��rw}j�VnrS�8͇��!�S,9�)Jj|�����n���������@v������$*t�$��ƴ�1��[��A�}	��2���K[JhؘC��:
���&K��P ÷A,�9��^	�O���fl�M�8�^ɦ�F�kѤ�!��ys��-��ψҔe��bׯ�n�9���?�w�c�"�XlxVHYEB    ea93    1880�����^��ZQ��=��̷���ڬ�sڴ��WU4аO�݊�=䲇l��⛟6c~��R�T%`xa�zv�^�M'&�Z����;~���%���w1�IJ�q�lc�C~�8��CW
���Y�1����_.ԝM֚�L�C�@�ro��]���ݵv��$ �$��>I��S�� w�عeT��-�$�'�������N���"��z�V��14I
4�5�@���hSzQ���[E��#�]���v+�B �X��3og���v��.��̜� 01�h�y�t�Bw�!�yC�@t��0�>C��kj���Pb�����Ac���0e�qe~1��)�V q֬� x�9������S�ME���%����K���`�aF$7mb�i���T�do$���/f��K����+��*��.țFQهC�P�i3���^�-rrrm�L@_��B��W�$X��}�O~�#���)d��*���q|`h�$D��MU#7���R���!=�կ�	���q��Ӝ3Rә	1�VFv�9���8&���(7�Q}�D+��vbU�4�x<0b����%�~�� ��!����v�*��t*�]�1���1^{-�f-��z���:� p+3��T�fc-UrA��?�ܡ=:���3����]����7T�Q��F��󊕲��V�Yhd��'�>��[F+ݬU�9���կ�*$O��dJv<)N�T}�H�p�[0'��R��3�zG�zx�{<)���Ʋ�$!A�r���� �j8��M�o�|���`�Z�L�߆ˣ��-UsC��
��.}E�����%���i���]!5�i� �����5�\y?�ג-t0DpS�{V��-tڵ��3�+�����uN�EVim�('|ɢ���(�\r��&�7��q"V�ʿ2B
�	�a�9�7+��F��%
�Y���rWC�B��,�>��Wm����>r��]� ����Юï�!G
�=�*�N��;���(� 0�������V�a��V�P?�/]
:�$C(o�P��r�06�9���
lEQJ���A�M`D��s%R6RbBm +����~��ѝ��")T����!����x�?4=9���|3G4"���Q�x����a[n$��s������,K�|:���
��A�� R��}��]XM%BМ���8?�xz.m�m�7�}�ǒk�?�P���
����2ؤBx�D����xc�{�:0��a�ɿ`.�>RTR��ޕ��?D:
�ލR�7��)�j�G��{1�=�F4<��6ٝd�ˢ#�q-)����!��'��Pt��X`D:A=��$���h-��B�8��o�XPT��Th4�;EyԖ�N��Hb���!��͊�ŭ	�OW��~j�]WI���v�����v�I^7j��
� �K��J~���5d���۫wkL+�롂 q��(7au�A�.,2��+'ɭy]���m��k��؋�*�f1<��Yz��24��>b{�����W��P9E>��'J6LkdWJ8#;����h�i�j���r�cZծ	Y6��#�h	��)�ڊ>!����/pJ�p�j���"���j������n��S8پ���ǂfv�f6K�ݥ��0P���RE;E�����Z��dj��-�o�}҇�[	,���[,G`�j�!����	ڐ�I"�aBﰯ�����=�;+%��`�*����V��o�h�0 �P�f`ob.N$s+�lk�6�)LK���Os����@ee�i]�P4�K��Č&���DͶPe��6D�S��%+�]K�N^�p���K�G�;h��C�M�xR��{pV5K�\>NgP����;~�����|P�j���i�(ܸ>��%���?o�ecq�y~���/%B����ӫK�Y��4�Ҥ	"WH`i���?{j+����D�%ڷ!Y��R�#���u{)��e)���f���~�z���Ψ������@$��跂D23��9� �� ?;�L�+b/S�l\Uc�|�y!
o�=u0e�T[��ǭ k��Z�]X;[[�ׯ[�Y.���Q���]�z*73 v�k����)�]
J�����~�7��zv�����A�3g1\b��n��R�_���]^�P4�ҹ�9����S��;W�B�$�� �h��pJ��b�Q��ή�?(QAs�����H:�m���I�\>���?ᮩ¸��9�y�|�B��sFKNHRj�ϫ`�%)�}���K�;��~�9<�3�D��e-�2d?��Nd�nc�}���|�H�,s�z��d:�x�Z�:1�i��D�l��B?+k�{R$0�E�ka���Q�1����'�c�W��A�����,;����jvF����"�%=4��a״Kσ
�+��k�of�Z]�K�\1����7	�A�܄4-8�Cӭ/(���rP9�������xF/�)>^X V\�rN��|�*��{Ӥ]�9^�e1n $���ww�y�㛅�{�V��y,ԑ�θ&2 U�7����I��qW�=�(P�~k�w(��c4��W
�¨�*�<!�<��Q�_e2�)�u�ϜTb���H�A��O�m6w|�c����B�L���s1�u�S��n��R�j��"�,��Y���AyH�嘑����'X��NşJ���ϊ�5��'�ݚ[�H���}N��L,(�XFԛ�EE�󝬻8�`*���m�iz�	�VW��z�V��j�	ʙ-����@�!o���8��'r��z��bԯs�!�D��Zv^En����i�]fa�p.A��&�)�T���Y����~R)�!�+h�4a����#�̢�3�#��e�j�ūy@r��O>
��aH���3a��Mi�6 Yx���${��')c
�U�	G]a���ȅ�w.0_=�ȵ��J �;O�#k�� 
c�i�%�{/a8��>�]d��Y�<e���P���Aƅ�c�,��<�6pwߥmW�1
��VT����	���Lk6���c�`��I: Z�K��4�[��H��
���%9@!IF������i�<!rn�	�I�	��K�-�>�����X%[��x��b�A�����N]����栒@hp�9Ζ}��I��\��� �/���Lyu|�R����gV�_�"�����{�b�I��%G�j��Q��n)tJ5�� 7A`�dx���	F�="�W��3��h�D�G����%饰f����r����{��i�
ugn4�Y��<��='Ig���7h�zZ����xs��U>����&�Z�ez�m�T��xZ`��Ў`��Ce�TpWf��x�î����LV����A�5ÍH��N��y�����TJ3
g�QPo�dA��������%�I!y�۞צUҙ��%�H�J�ّ�5]}̏�k�\��i�`K�x���cH�i��ps����'ӽ]���v��������EN����2��3;�;��$��P�{?X����[ƣl���#
N?ԯ* ��"ރ�J@���g�u>���^�u[�sS�}�_�H�u����p�A#��Q|!WWe H�^��L��W3#��7�tV�K�&�4�oe}!�*�x�P$��д�c�鲀���b+K����2�K¾v��ꋈoґ<CY��8�&��.����){�qv�_�|�Q�����6pn�sAcQ�l|B��S�k�|�F�@�`�]^�`�̍ݥ���a�!�)
A���t��]= ی�}�����i3�S��~�w�LT�8N۞=�������IA�E>J�Ɂe/��e���l�-�yC��|�@n�L�$���H[n����U����X��l�@�E=�bG�� ����K��>���(��J�΢�(�)D�3i����HGO+�}��2��q�Jo�֞�X�V`형�JL�^Q����wb�т6��]��t�m�@�nW-[�s��dl�1(�T�H6�6�=��?>�(K��u�Ql��?.���1�y�P$Q@�{�;�V��<��d1�N��q��1S���mSc�c�*�^�l��N�n��$�+��&������Մv �_X��(�%�c��(�{�&�T0B�N��/�9_>z*����_�r2���&&t'([�_�|v�D��$|�u�>��^��&YSoe��2t&�H���]14�!��`&��O�2�!:�Q*��V���U�=Qo�]�
�B���<���	�/
��a��*��*�Tc!'`e�g$eU��t�H��^ ����x�$������G��9�O�Q;��Y�j`Y�f{3�&�e��+��Y����o6N{��u��ྡb�V@A-r7�v��8�M�ƚ��}�Jd�z|�=�38��y��]2�Z���ZM��	�ϳL��{|�tn�Ԇ�xw�L~�h�Njr�4�N^�g�;.�P��s��j��W�V���Cʕ�ܒ��i�,v�-P3ḻ�-t�����;��[�{ۉ��wCo4�ސ�&<�Jǃ� ��T�&����[���ڑʞ��]/9ۓ�:+�	wVڇ�Z��M��ڮ�1���Ԛj`��E�73�3�K��B��K��$a��o���D�5o ir�@F��Ǫ�� �oݹ�����B�S���&��<�-1m}=�@�X�#�l��R|��5�NiߋE��\���������JkA)!!��!�UH���`����M��ߪ$d��;GN�������u�CV� �M�U �{ف��O0���}^M&^7��}�ߎ�!���{����*o0�({�`��!$`X�g����AA� ����r-��D�0[�	U�#�}�Ј��N��@���Ɛh����A���&�WsF��'ȣu��t�� N=���'e�]��)g�5{j���۽l_gQ�Bu����S]Rv��P�\���&B�9?��p}���@���a��wl'���}53Bw4�Ow�r��I׷�Cch��Rs�����P��e��kq��cp#��xf0Tt�H�x�mUe7�?�7�ŋ汸QԵ��k8$Ү7/mxpGϮ��|%S�vF�̆��d*C�(��2ab�qË"�S	ǚ����+��5��$�۸��ߘN~���ZriM�P�Wv˱${,y4�i@L�h�!`�]Նv�QA�(�U�y�yso��ڐx�Z ���mg ��0h?��.?�t���� ��r̰�K�ζW��EH�@�[訬����]�Q�����Z��9#�ʴȣf�oZ�],���Z���)�-NF�snA��6�(���fSxc���xa��f��}'7b0��rV�3\��B�I>��W`��ҙ�N�C�l��e�j��q(A ˛sNC3���7���aĶ�&�\��4͈Uf�l4|��{@�`�9�`�q~*�`C�XKm&(��IcN�/a}���.�R�"Ƨ�u|ɗA�Dk��� Ȼ����F��u'/�omHa;x0�`7�x��j�q\�h��/�*�o�0����W�604BMi�Z,,�ʪk}j8�}���Ο�XI䒉��d���x~�Ñ�f����fB��Ԥ��z�����K��F���X������GZ�b!���MC��:��xJHQ�۷����\M�� �����$�R�8�.X�Ç�z͈e�߀�������b�F��T�[hW���SW='��w�� ?oF��i�:#K���n62��8E��9�&�1H�4ݯ����9ɢ��1�7��.4�<�N�!�h���"h!�z:�����>/�W�t���gY�8A���*�V�0�d-j�_o��߬�e�V��=l L	�k��O��X�X���i�`��h�r�_S�d)���.�W�/�b5Ԋ�q��ra$r� �@յIq� �p�e�����m�����턔Xb��$㮅�,�u* _���5q��(�;������/�P_o�z \�X�н�,Z�Shp�Xh�5 y��_�^J�a���N�L�����P,��!�S1���ޣ�a1d�舻�<�kd@ߩ�ܪj&�Ѩ���z>V<��F�΃�:&U<�=M{V����P�ֺrx�F�V�_X�3aO�M�{8��@���s _?���ݖ�P�:Ԛ	;��F�ӔBT ��
ll��5��q��k�G��<�=?��M�um�������7K��+����U�������>�m&�Y1[