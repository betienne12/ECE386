XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0q촖�}��㋔�q�O,����a�����*kl:u�|~kRG����x<)�h�s�3�O&ڹ�����_q6D�#rX�Y�U����	�v�.)8(6y]�Θ�3e>�����sc�,�t�@h��w�'2xW�+����H�e�G,��P���v��k��
�FW4SZs9=�p~vk�O�܃��&�³HKo?�����&�F��k��M�S�y�e�����Pv�X�����Q�fn��?2*f$2V�!�t�2f�JJ�<�V��/��C��!��~W�B�y���ޫ����p'���VٱI�-�41���\&�J't-~Rm���,2o����8b:�(����j�xvy��.�X�w��ZO��[�����u�B��(E��D3����*|%����������bĔ~* ��Y}� �2+�ʂ�a�dv�^�u^�A날�fL��H�x��}��'&�z�/<�V��%ԚT+�2��Kv�&��!���^m�+�fzk�"���>��x��peo�#��l�`�K�F��{�UMS��z��9��L$!�B!0~��}L���?>h)d1� �{ ��UR�d�`��@���AH �c܌e�CQ4����)�ǆ������8vڻ'�2�7c8.�2�6����hE���q�%�7�C�dL%�xǆ9L������FŨ�NG�U �c�׶9��[�A���K��K�
ʝ:�xu ��9ԧQU�r��k��������3SXlxVHYEB    3504     cb0CN��;ۇ�hG�]mS����P�h l�\j/5�J�k?Gt�>�"��AQ�c�S�V�k�Q���K� ��U3��ק�dKGg���Fs��y#��'�+(���x���4�~���S��:��]ͷ͟�$%K͊�����1i��Ŕ~������+���SsC�Y�|a�Q�Ɨ���z��&��� �jC��,ۦ=�)P��Bh����I5X���t��dr4�0�p���4�S}Q��v��K$���9;�#�O�Q�����h�K=}�y�Ŏ#r�ڨfrd+,V�R�{�2��ե�~�螸2�9�������Zs���� �j;p�Kx�]�Q�A��P<����NZ��#��{�"d�ѕ+1�"Р�)}9-��$�1�K�]����a�9�/ŉ���:_��0Eb;%�|X�~����6����3�B�>2ռ���$���G���@<������f�q]�j�����ܳ�Gꕿ�F�MsJ.	*#̘�sƄx��(�r��ś}.���O�����d�������E�#4���
&��\nο͖�E_lky�v+�~u�S���,A�Z#������;�m)�
�7�o��i'I57�[�$��a�,�����d1�=�*·�;SmҠ)��2��s�p)��`�z��M�A�c=U^�z�U���c�?S�$�h��`[?��DZ�Q��{�i��%6�CuTj�畆�����oQ�������Si���B�,�{wD7?�<yV(F6��q|����e�Mu,���Vi��l+�cȼ�>�F��Q��F�]���(ߜ���9E�;��Ր4cDa�@�����K��Q�$��v���2�e���Ը��������>��C� V���#I6[ܮ�;�p��&9G�j3����s�;��B?~�v:jJ�E�c}dkjl���W�=jl��&�{�5v�e�(%L���c�W�v�5�R)�(��l���ʧՍT���>b}�2y�p��{�
����V�J]���j�~%x1f��UA:�g@��́� K�Y�M��k(�TS��NJ�C�4�Za<ERWq���(O�Hj�^;l�F����[xha7���Xr�%���l�,;=��������&�G�9~{f��RR"�Zկ�q�lt���DmCZK��M,���s��3�`���W#����en�+-��Q���tqB��'w� �|�$�:�ur�E��?�2��9��3KDMƉ�3I�=�C�:jb0τO����E �H�|E�_P'��&G|(50�b9���k/������tS�J�/턻BAҕ��m`�K��uaJ+�%��S:���=�8:�}>�ğ�$�Z,;v��%�b�*;E��;��v�V�,<@j2E'ER"i��Rժ��@�ܯV��?�Yq���,A�+%s���dZ���y�����KϤO��~
�%�7�+�{\(��j����u��Jݵ�=���5�:E�k-������/a�Һn��W�9e��~�$,-��-;M�BSң��
�%�(m��3����e�,]S�V��&����+�t��x��%1��u�Y�1v��`��au�[.�5<���vY�R�n�I�Y)�f��Ǚ��Z�n��-��\�`pu/��&0��c;>H�.4q��ǈ0Q;��n?�e6c����0�s�,ܼC���/6̸�4�7��
�ǭ)a.���<��'�LS����#{ Т���v�BU�rX�B����-Jq�_�����6����h�)0ḵͼJ���F�����pC�?\HNl���!�IK��3�	����i���ЬK�O�َ-|��T�������������9R���?c�P��M�rnp�J�tG����TVz����lŤb �N�@�<�#TҒ��KK=M�ɿn�)P9��c��bӋ�FH��#���W�e��j���!Ցk����\�ʖ����r����K��Lɚ���j�p�[)u%���s�(��boײ�����>�W��hѭ� �[h5���(�})Ҽ���&:�r�$�4��[�I�a�0��L ���M_A�h�Q�pp�R���S�Ƃ8���H7�f�U)g�A+m��1��g�3�X`Hj�MG�s�-�F�>9���K��Ǯ?��s� �wf@#�Г�F��ǚy}��Ϲi�t��h=Х�3��7��f���G��CT�m�>������e5R���"���V2�Hr���(珧�r�X�Z
A^N��g��J.�rZ㏮��gg��-H�]�8 �!�D�e��J�>~d��p���*���~��ڠv����Ė�Yyq1��6�E)�S�H@�~�q=K�1F�qTۥ��Ф�VB�0ې
O�<a3ÈS��]���=��~�j��3iK�[?4J ����d�N��t��&�m,ێ���m���"�[�i�N��`�bD<�,]�2���Ì3���w#Ei��L�<�1�l������N4���0�-��",f@�����¡�4bf P�%��tN�In������t�H��4�\/�v�4ǌ�������$��( ��~?�-�\�|���iP��jZ�����E�d�jm�PL��P���|��U�N���~r=�P'��ۈ&x�ݹkjA�~&������2��Zwn_oS�~݅�P�F�([���=	�f]���?8b��#G�Dl�uf�L	K�����uΆ��h���Z#�4�Z�{�"�cs�l`�z4S�@��$�/�����n���b��l\e���-��N('c*�� �Jz���u����ۓ��Y���GWr�ğ�a�/�g�M�%��'2�@m��2].��h����@���j��+2���!��I��^�0N�^w@��&�HS�]=j>y�ܿ���Ulc#����,��gg�R���S0�M��0'���t�pp�6C�l��6&t?��"���x�z{;-\��f~}����-��w���jh6����Ա��(���T��a�ÌRQ�L�����<�sx��-wF��g�M������Ivd��|C¢�a��0|0̈����N�U|���Sc8��~�OV��(%�"uۡf�A���Z�ǽK(;ِ���b8�z�Q��sX���fY������k��Ӯ/.����ž5:O���!ޭj�hP�����6]Y�aP��-T�����W�r�_En�jn�?:�G���?T�q�A���