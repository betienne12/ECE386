XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����?*��ܫ#��W���ĕrZ����2����O(KP�^
ٳ#LÜ݅*�#y�����`�Z�� �AOT�(I��nVɕ���_���>��s���~���$� ܮ�?�Wˇ�ݴ0�z�MnO%.*�Ex����b�W��0e/ZQ4ꢃ�w>���eR3��=��<����f�8����̔!H@���-p������'�Ȧl���q�$�f ����w�5���,?�W;��r ă��>l��&2D��d=�Xf�j�2U)�4���� �В+�O{��
GOEe�f�יV2Iy��X^�}q������V�Kp�T�X3�oٝl�	�����{1��;���M� r<�QV.sh��OI��� ��YQj�)����Ѧ5]Y��/�^<��Γ{��Hӡ�)�]����5h���n7ya��+�B��e:e1#.�(l@��� ^��Ґ*a��--�UΕ��DC����b��//)�0V�ѫ��DZ�T�b�Q�4���N�],�B���$R�� �f%�xJ�Ϊ�c��Bp�8-���*v ���Ƈ�Є�.s5�4E��"���V�5�ܹ���c�3PDW���������AiZ$"ŵS�����%1���E�sb��ZT?�^:s�8�� ;8���W���+e�:�.}ٿ�JAF�ǩ��W��W��k?L�P?\�n-�_�����<�(�i���́W�6��p4��.2qrz(�r�z��8�~���bXlxVHYEB    fa00    28c07!p�{��yL���h�v+#���*�I�q�*ԁz�^��v�&	_�Q6���N�����a��V��G�F]f\8�����1��_i�ݒ�Q=ܮmv��d��e�g��|x��x&���6��'H<�-7��J��~>+�k��]jP�w7ʚL�B���d��7����&����I3O����O�ԯ�sBw֣��{�m�oV�?�|�o�ؓ6݌u=�Y�6��������-�e�
�|�+�XiN�.����"9ޗU jM;�=�fM���٣��GR^,8<#�\�3U�N���h5]���W(�k"���ѱis�2.�8��z:��r�G��]2h��	Z�
X�d��hM�Ĉ��A@~���_�}���G��. �o݌::PU����IJ�7��O͊�5��5��
z/H��g�a┱�p�l�7BN��7���B��7��,�nG^�c��.��/Hz�ELR�&nBf��|!�T�Er���G���Ñ!����N|�������\��L࠯�t��7dn;T�<����n�G�y=�6�z��:Lp�=;�D�!WЭ~X.���,ʔo�ԇ���dZ쿆I�V�фv-�.����t�$�x�!��A�rTT&��0�ݣ�dT�ugPX�Yu�c\�{+ۚW�?d>�!v�s��1,6��7��+�lOKu����8�˸q�9uUt��O)���b�:S��Pr��eU4A�v�Ӿ���a���PD�$ �1W�.J����-?���͈� E9١|���mg�Ӄ���)d�P�L�BZ��8,
���#��l�y�b�$�(�-�p������m���y�{$]�nJ"6k�l�"*��c�����'���p�ce�Л����B8t��諣�zF_���U�׷E�Y�B2���Р�b/5$��* �A��8)�m�E�x�9%~��;��1�0�XtMB�jy���.?���P��t�'��Z��ntC>
rG=�� 1mg������oL����/{���O<:ɪ�z��[��MNQVM��JB�|B�a�*���QN���(㢚�v�8wU�hz��y^m�%rc<Jb��_�%2�VO��?d�8xk%���kp]^u^[��-��3�cY��o�[R���϶'F��U�R��HH#��ͦ�[	,
k6ϫ�˗�0%�3�V����>�&�����N�%!��E�˷UbQ� ���4�q2���5�Z�>b�b��ڡ^
}4��+C�p�Տ�Np�~�Z�oq��4x{n�w�L�/�Na����u�r{�ʕ�
���$��h~P�[[�o�a�HЋd9�4�s�X���{Ƚ7櫲�O�g�%dAJ�V����p�J.�VZ7����fs�����z1�ڝ�N��況Pّrzp��L�H�[Q�?��^~ј7U�𜌒�ݾ��M�fU�f�-L�~�}��\��btU�p�^D_��`�~@��'17�L��Z��H��q�x�|�MM�Jn����F�����vgax��K7O[d��'�R�M+��S
�2�
??8n:R�x�ǻ^��q>�C�{2�/��~�
|���΂�ΰ�4�� ��]C\���$�%��X6�n�qrB��,�nj�1���#f6�t���v�8Sɓ��7�f~X���u��A�k�6�\`�p�{V����!�f�M����x�֭?S�E�~��{��|ۼ��gX�e�>�z���g���0��j<�i.������i>�(SL�"h��ߋ��~Ɍ��X�����Q�rF]�W�/�|v5Ęl%K�s�����Eɓ��n�N����n�6K-�뺽�0v	U��0��?�Ri#yiG��J���+�͠A>��R�c(fca3HL`��5p,��10C�� _�8�~���8Fmb�����a���J�pmy:��*�Zpz]F�G�d&���ܝ�K.ŀ�Mo�9��F >s�ێ+�gYEN�2S�6�aL���A?�^^Պ<��s_�@��DL>=�Ύ���֩P�w=�h�ȳ�P8%�!��b~+s��W�ׂ��Ũ���-�W!�-���n(I�~�aڠ^](�w������J���� ߅;H��.�G��}ZI5�N�R@�p�@����E��2����6ͩ��2�Nj^˟� ���*���55�ltc	�w��g���Dn��B�4�6!ON�7�%	d-�#*��*�C
�7>WbwP�W[aWT	 P�A��D4�j��wY%���?��u�Y�KG���$PS����8��J��{�q��? D�1���vy�4�#z*�S/8�cf75|)�9i�o7�ʼ�.;l#o+"���k���̀0�;�~&�p�K����*�d�Ø�%��z�q^�sˤ[��.0A��}��YT����Lm��H������麐�
V�4��;:��>:��:u&�����5�~�jg���k���,��j጑�]B*���nj	�qfV�#W �x��l���L��P͵����U��D��-����O1$3�E��r��a���.���(J3�I�k*NЅ���K��{��Ù�۷���&���~b� ��)^J���F�����-Z:5emԽ`�PiҨ1@C�4@B"NoM�IX^����������u�N��KΌ� (�2Y@��b�� ��Uj��X��N��5��	��H��v���Q���@4�g��~xYrȸ�~&���Ơ�(c �M�����+��/�O_e��aٹ;{������$?���2#pؙ��9�,N/V2\�X�omhH夗nI����p��3�������^XE-;��w�/�x�)_���-Ȧ���n�	C`�i��$�]�1!�t��5�B���䲫X򔤟H�DF!��� ���-Uw���
2�̰E�&�п�Pv�xµ��-TO�v�՜鶬#�
�H�D,��q���#)-}�����	��Hên�D�On/R�J��o�\���'��E�L�5�u���2e�ňṃ��К�"<�Cx���
����>�U�y*ݞ�#>r�Ȕh+K�e�O�-��WB����go��m&�Jפb�E,z���q�Z���#���V�}b��2F�$���=�ӕ> g���n��ڿ%�����]����L)D@V ��pV1{�d�L�y"^#�	Y�� ߷�>��3�':������"L�e,5m��w��B�a�+�BRYP7 1����r�?�:��6~|@��k}1Cׂbx����sR/���vl�0���i��VK�1��2�p��^^�fg?��7����w(��˓s����u=��=$}�-)�r�V*m�� $ߔ�h��T������Aԇ��n,������@WH�Ѧ����u'gh�s�2ʞ=��#�7�ｷ]V���i~��	�X#Z�+eğw���F����쫯8��,�>ٶ���!
�b�J|Ѭ3�R��C��}���.��7s�-(�Z!�����bz�U+�+��P���$��.^�v	�*8N�]�|$G�K���#�3孚u:έ���Ҥ3�u�H`{*�.��f6{O�/�y���A
 �qտ��j�qM��B)#����dbD�fOm�I����F�;���\�Ŋ�,��1�mw��S�{�A��ǫ��Ӳ�+�0�ۃu��R}bMTs�.�.a>�����n<�t�V�=-T����v��X~�d���e_r�!������ڌHBLa�[BD��|��Ə���a��
&�a�I�zYsCy��2�vً�F>a��l���]��f����iC�����K,�ް�p9mQo���7:��̵*Ȁy�&�䎶��X���7	d��&��DDI3浟l�X�ըE $*ۻ���ք�i4�8zM�nE�H��1�bd�0�	�b �-��W��&��N�_{V}�?o4\_e>meB����j��� |�0�r��6j�lq���/�)�^��A�/�[�14�]�g��b���z3�����Sى�~A�p+��I�b1�R8��;:)�����R34�b�B��fL�c�V-v�]`U�
IMA�k���ş�l�3+���ע^���5���'g0��Us��'=�c�A��MYJ{xOt_Pc��{�AxV8b�x��R�h+��p�g@
9��[��һ}�j�񁑻�����G�R��������| L�yi]|�pR/�nH�De��%�Q�U3�~|�	��!~<IZM𒨥�8�!.�
π+�O������~������c�E!�/�C�O�4�����`��S�P?�_c�{�u�#�`�ɬ�=ې[���3�a��c������1JʟR%1�� ��	cT��*Kp��;YI����5�<���V~l��� ~E��ޓ�����#s�QʟfͅU�h}�K���p�p5���R?1�y����V�y{�z��C���p�A/��ማ���w�I��ى�������w�7�"�y�4��0���}עg�l�����/A���6v�]M]�Ÿ��F�#�:N�!6���$P���Qm�*�w7|����-s!��uУ#o���5��p�x����� Kr=h������}��fK�B�m�F��r�4�,_]��ͭ�֨�����ȻGJ� :³:v�3j�p��K��D�n��qE0��p�{�Kā�E��� ��T�؁��1?�\�v��p�ȁ�/�֨}e��j5pU�k�`�_���vvy�s�m6i�!>�lT��x�C��ɰ���7�#o[�-AU=�z���� �G3"��������	3�}&�����CCvs�A�)J��m��V�|g����˿m�H*w����l�މ�A�F�2�m��.%�JoOi��Gj�\��f���5�����Q��8�7^�$~��Hh��#Q&�끩+D���qƦ���Iv���`A��:qY�uX/��a&��	�춼Un�f��ȗQ?�+l���{� �EWV�;���:���Q*�����/�o���7VC�Ȫ0�Z��Q#�� ş�A4�����)A� �r�qd�Q..����y�w�W��s���m�M�ep�0G�)��� ���9Ma�ݟ�L˃=ZuCj�l��o	.���J�Uy�8s�g��	�~�M�˟��$�@�3$J��==UZ�~�%���Bt%����dU�8pq�X�p ���k߿g��@��a�? 'TS�ѿc:�d��mo�u�@?3� ��}C���
~����Η
"�3�wP"Z�H&�>kt������0��J�E�*o�ʓ�N%a(��#�搹<p�6�)|zݑ�L�v��}��d[�������Ppj��׀��m�F��<{`G�d�h�����˭3}\�8!&��-�����	����GD��Q*��I�xCo8����S̆��O�¡�g'㸢v-��,���L�A���ze/~$얁;I�KF\��4,8L�ү��S�����FZ�NO1��ۣ�f��9�6��	��'wv�q��4%�k�[2I�$��o����*��8n���+�"y��_A� �<nŎ��MGCܹIm��)�[l/�G�l�`�n1^�}rI��iA����k������������*��t��O��$�GD9�Յb/,�C��˳
8����;oAH?榰��Y�|]�֓�H@��=��W%��/�e������q1�)�$뿢L}�m�Qݘ���g�U�pNG�(_�凶`Bn����^��YY�E��#�Aym�ӕl-���q���PK�}
����aM�K�E`�b��x�i�^�g�$�у~�J�M;c��aGW�U¦S�w�+�����oF�b�������s� ��\���#��H1�Z�ڌЕ�)4�k}Z�η�答�A�ur��,%��m`���v9xr�+R^������ҵ��[wӹ��F)�����W�����~����?�#7��+��D����Ǟ�(@��ŝ����j�q@9�Y���f���ʬ����<����S�OlgӊE����`D�%���'�p}e���޴�S���+9xY,���8\(��:��G��������>��+v��BLs)��ŐI�S8ڠ�G��~[x��Mvf��ȕ�2'G�����ͳ�����h� ��\�C
G�) ���	>�Rč��-��ռ^vwi�_��,��&\�M�9�>�;���i��A4q�8��8J��Zn-��I��ت�T��Rni��l��0�u~���3��]:�h�	Af�	�C=�F�e�Kp}t�Q��(�+]�i��}_�u �~��|B���=Q�N���Ձt�`���o�e��������֙[���|�簵6�4;�@�����Z?�_+Q�}��$�r�A��kF2|���I�\
��ݣ;s=���G
gѠ�A�3����(��<.�e�B;=v��Fa^=�|l� �C���;��G��اD]�>w�_u�TK#.�k��Ϟ2���X�	ľP��t�\Ml�K�D��c}5�`�<���P���
4c�ik?H\������V��W	Zld^`��\x�{�ٺm����W|�����_[*Ȗ�ε�vvM���n��Le������Rd�{��9����U�C8[;��${hi�-��,�����M���Z|0� Hn����i�)���L3a�t�{�L�t�\5ѠD�J>�H��X�,. }ļ�BB�Cd��֡!�<����|!t�t�����3-��ҡ�OD��aI���$��X�з��M��T
E�"���������31� �4 &��7���P�&���G�m�ɖ� �e���r�]ӌ�*��+��kZ�^�k�8�&�n��'����|��A
��,�6k�plVh4q3XK/�L�#d�������ėh�|O#R5���{`Ag�η��K!o�R䌇�ҨE���B��ɇ������=0=�N n�����(��M���)K��H:c��c������M�Vf=�粒��Q'F�=��"�õ��~�^Y�� �,�kF��*�e���Tt�{�M1�_����.�	n'�n��Q��U�2D��i�oH=� y�c�s/8���X5��x��U�ϟ�����,�E��I��v,��t�܎�D��1�c?�Z@:z�Z=� W43C�A �	*\�����3���Q��W�ɉ�N1s�{�),?�T��_[����m�����!F�j����~PO�_�ϭ� 	�v\�յ��E���G�[;җ��D�[��,�G]d;bw=l-��-6�Gl���2đ��JK�6��:�sN��<F��Ւ���Ba�}���(�$�U��~�3��>�` ���G	�V��JJ�����ك�$�ݗR����N�Q��lc%%�#�~�NM��	��g���mC��Bt��&��A���\���;ڬ������O,p/Q�;t�����-"Um
���Ī�i���:�B���z`_	��ؒ
��w�"Z{(dDoUBB�*�A>x[`k��R��A���0Aܽ����<bp��Yڃ3�٪�bγ/�#�2[|�����e<H\_v
Ŭ�v�[�������U��{��t�C@v��f,qf K�/q�7�<}U#@�kD�@|J��v�`6y�-黤K��eY�Ov�׿j<F�u��cm�8+�N��o�i��Wt�F5�<��g2�tk.����i��ǚf'��9�b1�L}D�܅�a���t٨{��8�N�D.�w�9���
p�M�S�� ԛ&u� z{�9 ��e#g���R��!��8�ύ�vѣ�bx�1�
�Z�C^�zSk���ң�o)�%�����f�4�ޞP��0#�R�-���U�h�qW��o"�&�)�K�ֶDA�^`,����m=�ZW��C�\����!�5o�̮ k,tQ^�s�	D���.ݨڒ�ɥ��2�w�Xn����_��k�_��ـ�r��9~-�������X�Y���lĽ�h��RxG���u��%A�F��RB�x�����,�F��,�V\Qݳ���r������r��"1;*���^o���_æ6D���⺘4�%~��J�UK/���tV_:}��`m�y�׫����c���F\ޅ���32�$HnV���˗�hʇ1:�j��� _��;����-r[9I5v�Bպ��>D@Q�o��cK�gr) qM��pt��0�I��vY=q��aӴ��=`c��������0��v���U�/�cI��>�X?�8��#-RagDy�Jo!�&�Ƣ�r�ю���s��H+:Z���$���U%���{�F��ޮFt�^y�I�˄�+�Sَ�'fIz"� ɳ�ԉ�G���m@����@�+;�9I��6��Y3��-��j��:�[��˓`{Am2�(ɂ����f�F�L����F�.�?%��{��:��x2�]�p�!C)ꋗ���%�J����R4\����5�Ta����҅1Ե&����mڨ��)��*�7ˇLxD���ES7�G}U_���y�1"tn���$l��bT�*��I�e:�4GɃi�/�2�~)�ya���u}bi	��Fn�*�Oa��܌����uvz;|0���&n�-ؗְ�{���?w�~�c�ƅE;��е�Kv��qY�(=��9�إ���x4(+���IM�=��2mH3�;$�px�pl�cy��}�8�E�e~�EXv�Af}�fV�����޿>�~� �N���F��'��=�U��8K���bl�S���>� �dP3�g������kPV���Sf���.,��k7�ȼ;���G\�~��`�9��a52��@�|Zd����Z��9*a����ŗ��M�+I{����t���n&����9��w���O�wg�SI�jqv���9 �(���@�[i��|�1s��*������d9��к�.�������d��z�4��ք9��lp�ӝBηk�q�eܐÿt����M�{�����;jҵ���U����"\�O�ŵ=4��7��Im1��C�)ح�������Y6�h�P�hc����Ĵoy��i����*@$���y���qO��k��53�S�٢�3�����r`]�����E�u�Y{v�m14����
2.��寗�O�%��o)�5���L�xR��9d�f]K��d
F�D�A`�R�ix3�ޥ�qà�?}�h?Y�%�7"�7���i���2�w�����r�O"�+���ww��ܳ����@c:���fI���7m�^Et�	�l�&��_6�GnNH.�8��}�	$éY�*�$uRH��j-��W�g/��Q�[s�k?y��C�,_�4��0<FB�/�ECJ��@I6�*����3��P���J:� e�k|���V)\�@L���ߒ������Gjڇ��:?����L���WR01+�����焠�W\W<�$��C��v����8��		o͂aS����a��C��~-�~���� $S�,��KW�z�nb�!�=�D�e�^u$��덴N"}ŏ+)�92�D��-��D���w�E��b�"Cb��u͌��9(���3T�����V0�m�b���Aڕ�q@�O ���)�<1խ�O��2f��>��,��Ȝ00G0_�*BG �;��q��(�����3����W7���v�����ǅ*�O<\ӥ�Dt��2	N�/��Nq��:6����2��U�]$S,w��C8m�Oꓩ�@+;��-��,vo&r�8����_I��TO9����'��ĽQ5V"+&!ٸ�n�f��/�ڕ/�|����D$ -*���
����צ�｣�K8^�	{١�����yf�8$�a��Zp{+�Cy[�k�TgZ8Ѡ�G`rY���10D�^բ�G=�o�R��rZni{ Mٓ�)���|2��C�dw��7�ƹy�������f��Ra������bG�CMɱ96�J��9m	�ިq'g,2I��X���f��~�g��jţ��)	hpm`gC���:./G��Z�_)��?i�#v be=P3�r_��S����.� ��ufv�ɲ$���Q
0����][ݛ7|���/����yu!��v ��x������J\��]̅������Ɣ�)۟��IjD�]�:��Y`v߸��0�%�a��5AO^D�>�C���{������/�}	�����V��[���3����tB�ѧ)m� ��#;�Hrn�Ċ��D��)�����C�]2l��Đ��d��s�!/^[6pH�ua�/��~�O���V遝�+�)��-_:�I;vX5+M:����ҁ��	����r��Ѐ"(�5l��ݡ��0;����JXlxVHYEB     896     280E�1�)��bbC�|���DDD�C����0����bX�m�q~�
S+��l�ƮgiCu��#·��"v�ܕ�~�#1����:��"�7G��(iVy��v��˭_ rImt��� --8U�����DF;X��?����# ����U6"%�W/�v�7C� ^�_zl���/��+�#�-
6ʧ�($������)�K��F.&̜U(t����ƫrB��7)E/P+lk̓�2uJ�ך{�ïs�ԓ��!��=^ye"Ͳ�lI3V���3Q����f��=�Xx �蒵�_p� !�d�E��;J�6rBA�
��n�	���@���;���%��" �ʩm��yFf�=/	Q���ۉ��Z��{n����Z�s��?�@/��^V��]�մ�O�Q�a�����~@�I�N��>�_[a+��$6��{��Q�O�:�����% �&K��ǰ��
0���E�v���QH��1��F�փ�ѻm{�X8�}�ݧsc��f���jՏ-��1g���>v�*��#�fs���/�B9�魛=�o÷ٝ��?S$����<��8��h���N�k��vN���0�e(���rX�υ��+�્�,ل�%��1@{ ��u������J