XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'��f8^�P!����A��G�1����&1L5�7w� =���r�n�xڅZT�[��U��J[ĕ�f�X}��5�%N�z�zٸ1,VDl;3U��A7�/%�e��*}k�����${<=\-�&��Wd�CX �K8�~Fr'{)/�t:"@�Fȑ"�P+�c�=����;/^ݒX`��*���AF��D�(����pV��q�Jר�� w^�5��3�E���>!X�2���Ld�)��b�A7�WK���j���M�D����Kԯ����Rш�q�4ů��Y�)G���je��'d�P�yֹł�������{~Z�����ṳ��*װ��6w$TJ��zT+�OX1\��=�\�"g-[��Ն7>�Ӂ���\������-�'� �.�f�ba�vG��V���F�u�w����Ŀ���۱��]Aa[���E\@^�r��dm�� m�I���V�/ӣK�~{�S���"mBo�E�!^�O�rHh��!���A�T~���� ��g���جQ"/��z�u@�ߓ�[��55�2��#��8��w�f'�h��Rؘ�i���*����&��4(��*��ҥ����Z��>�gߐ<AX�B�=pB�g%�HG�4��%�)jP���"Nw�����*�<U��*(�czO /<>S���)�3��v��$+B��v�FV�z�.@h���� �N7������5���Y�"&�oUR��0̮�����kE'�i����R<�͠�����_kXlxVHYEB    fa00    2260d�w��)��I$Z�.u�S�/ �;�����*�Y↺�0zP�v[�av���u�ǜC5ߦ��xI��2��J�8��9ZC�*�So��2
`˯��s���s[���c��:��*��X��q2��<wX�>Z�Y�r���U.�E��P��_�=��(�H���R��uƅ0�(�.�� Ke�o��{ͽ	�\ 3y �.��p�P�Y$�:ػ#�l�
a���tB\w3��,$�`��}A|�����:��ߋ���m������\������0��]��v��`3�.3:{2:w}-���i��5+&�qtMo����_�7q�l�q�Ͻ�\�5V���A�#=ru��I�kl�frNX8���>�-eZ�Sx���iG����a�hLЗ���t����^��u������4;�$����6�$�4���#/D�ӿw�A���N�[X�e�TM�>Y��,T1(P�-�B��L����T��fB��,��5�*=�e��*�AT��@��NS���tgH������>U�����F���֍n(�m�ea*�;9^Q�����L8Ѱ�^�~�g�dX�NR��ɘ��m�j$�I������/y�گVu����^�>u���3��^�Ab�Le��ڼA3�a�_ջ��<��7E�K�y=A���԰��_���Tm�	e-���J<�y͞+��~6���"(�BDw����;,� �E�²T��ik-��8��Ó���0���*�A���<c�E�r;�c 	��̺=q�D&kx=A�|�6�;Y	 +�K�э3�--��M��ڌǣ_k��#ō����U��]�2hm�U��f����#�AD�H:�R�5���>8�%��D����Oԟ�"b�م���ih�M��Ww�v�jر�y���!�=����ȴ9jw	�ڵ�&�qu�ޯ���
����"�(�W`�WZ:�շ~���X�E�ut`�PiJy����M�����7=L �$��w�ŒDg��t�9�@���R��S�6k�8�o<���J���	λPx#�`w���i�5|s�����R��n��!�� Fs5��F�E7{!�� ��<,8ϩj/��kW�a2��_�Yy�z�r�8��~��S��9Y��R	� �-��v�h��6���Ȣ;���@��g]|	<��VK��.��?qx*�:��_�[�&�&������X�������+y��>E�>�	`,��|	Ou,�N�m	6a�iPQ�O��+W���q��w�����@��l[ݹń� &�ģ16�.��F��A�d����-�Yv�����s���%y��@3��Y�!A�
���T��R��㚄�3���&�\�Ƙ`��d�M�Q!g��쇍��:�,Uޠ�s�C;�Sa7 ����c-����M��L��i�kM�e "�{s����-�8/�r#�z�U�"γ�`�%�f��"��B�$g��	��#� }���M�C�Z�0R�jhqy¡��zz�]!�p�����%�H�����D��ӛb�A��MH-�����}�;3.�mF7�A������n��/rd\`J��9��NP�Y~؊<��)fPA�Sד��^-�玻ku���4��g'I���_�,$=���$�Q�Æ�#���qV��Ž0��h�(�d�И��r�m~�Q-5fd���'����c�AbB��Wj����
�{xs��ǥ���>�u�N���# ��nj/�g��z�h�x?�W�*!>�b($в9՟�^~d�$�V�n	)�[��=�6n����x�*$�N\)vɰC_��U�66������$ᦔ3|T�U�}�P��3�d�%��'�4_zB�c8�1{zSw�;�R
��H���`�M�dP졢�S㖙B���+�Q�������{����7��j�yg�Xݏ�B��!���7*�%I@N���$K#���X� �n������E��7�l��W���;�mK4́��ŀ�z�BT�@��5��o|������9�[�5�/`�ԁpr�����J�����o�SXQ�~�[Y�&�����ބ����Q+��0V��#��U�~�]��)��QG��������eZ�����~��H�G[�`KW��Z�i��E	1w�Mz1\�S���S�����T�B$
��p�-����VU �(>�]�{��u�y��[!����b�~ %j��Aw���S7��=*g-ޢ�'}��m 0�����<�z�+�<4�����,�J�s"E-���oG���)��^�@��s_-W�Ҿw�:i��t�,�:��Q��J��I*��wN��~���}�Qz|�j��d�y�Ԭ>;�s睆b���Z�,.��՛� �����HoR���E^'�H�Ĭ��` �q�����Vc��k}��Y�-R��$Μ$B�{���;�T�H��Q��ى�n�G{i�^���,�¢lLM���I�T$+�/,��g���o���so���6�������� ^�6 �]�n�-3<D�ն�� ��vn4U�j�������B�z�ŉj~��
�b;�sjfF|-M�j��X2HvȦt�q@Hs�{�V�&0ʓ'��gcq���NU8)�k%+!��m���	ts�ft�PR?��B�x�v�$T�r,(-�#�/&>���(V`{�F�ԙdha-[^hU�����dш�TF@�9�N�[���L�#�7����,�N[�3���VHMj!�<"���œY<NcCzČ ��ooɃy3��2+ܘ��P�'4�=:P��QKv���e2�[������@6��uO�����	�^Z�<� !�����~��o������V�0��~6u!+��^�喺�;�h{̍��	)^*5~�6v���O|~n� ݟ���s���t��[(0��(�vs���K��C�8#QK��=&������l��g�� }�JȾ?�xs�{�/-]�e�$^'vd�`x�f��@�v��1�MVhͽ���-�|�6�VhL�La��[��6��'6a��ex��$�H�j4���pd�;�}�Y�1,��#�T�� ���~0w�a𩎪�Z< wH��|��*��rҌ3ήu�A[ހ����^/�f�V�rg�;���z��� �BR0R�b�UJ6��a'Ӹћ�g��^jݦ�h�V�:'� q�4[O�rS�eo��uq��0f�*R+���_��6W�{7DN�_� s)�ԥ�4�bw)/�2�E�9���Y�?$��r�EH<��6y�f�9x�|�����F�>�D}�1F�߿on\k\v��zA�W-��C��7Y���E��͋��C'Ͳ��&8��PQ����k��9.c
�HU9iI~�����*Q��S>M$8o�寰:���7��[�+x(P���ͤ��}#|8X��2�|Z��ے԰R���c����FC�̢�\V�B_�ezX��q��/�J�������2 �r���ś��4?M�(�?uJ�D������#Ze��.���,[2Cf���{2</A�R�]����p=c����4�������Ui��U^?��CTB[W�`Ӟ��*��#����0�/��J�����������h�v�v��-�e�� ��<r�(�\�,� �g�O�}�8\f����h�J��8I�w���{�O� u�X�T�{t��Y�%4����N�x���H�@U)�R���v�D)�v ͡]/ �H���x����Yr�F^A����ғ�}�ѝ�,c���:�эr�΅)��(��@���,���-O�E��g*D�#/��]�U�C����g��� ؃tVN���?!�ƈ��q����s=
�B�gD��뱡���m�E�2�?ܝD�@IG���h$��L!�Q����6��ğ��Ӊd��2���F�+i��k��'S��{�(�#��Z��kHf��R���i��ElK(3��V5/K8�AYq.��&֫@o5�4_�@�qZ�|8%��C�.�g�J7�|+2Gِa��� �z��M�-3#W�	Dni�'� �s�á�`�� ���Wogvl�T��t�u��Q���$�=c7I�ἼϢ��Z�xbp��|%�r��,|�z#� H�C��P�����T�A)�qٝ/�N��tI�C?����<�%x��tVk��'1��9���۰m��Yu�'���/en՜��e�Ml��E�0D	�����4���Dg��a�������0@zp��|R��֫��E�8��C������o�}#�"��Pf���iq��G��U�N����X̖��,��^mF��bw'5�R�&���5��+ �`͗���n����\�2��m������-db;��;`J�T��N�s����G�hBS}38��1V���[V��	�\�Q��J�"�%�ؖ2�9\�<U3�����e��(2�0+=�4�Єؕ|�y�;��hrx�y�ы�N��{>�C�X�nk�r�'V�l�|7�)��ǋ��L���)U�aN��֋`�ä)�-��W�wQA ������[R��Fղ�ﺿ\�B��P�rl��D�%��x\G����dK�5���A�:q�Ԣ_�$��Wp(H��:�~��dldS)VAs��8{Q3�|�	��H���\�Z(2
Y�)P�$�c���|���[Q��Gs�}ݡ��}�RИ1wBjH�k{�����0�/̍�݆HoS�m��f^�X#�߸g�% s�V8�q��@�x�)RXa�'�9�fY2�X�2c��ޥc�ء�֩�M8R�~���V�y
�� ��ek���f
�rG��^��5�����R�Б~�@��܏�]��S&��k���^�FAL^M�G+I����4A�I��L�A�>D�AS�O{N0��=��,��I�TW<(�V�*�w�I��/ူ���ƫ�lqϛA�\�YxV�n���#��I����2E/�|$�b��r��	>@���}C6����'2qi���8��ˋO�0}"�O���`�[������
�ZD ��>�'&7ߜ���|Ӑ�H���f/��z}ߝ�,�[&^$���w�5�S��8*)W���6���>����"�n��mtZc��ӆ�V��q���V�i�
<u���t?�b�����}!��� ������IRRӵ��.��'��B�@dj1�E�1�.+o�0���)
 �>�d|��fbNj��Ď��PZ�I�!+7=�_ɟ:w��l�����6�/L�N2�Rr$k�a)kn{ @�.A�#gng�B���\�8�~�"��9X�-�ﭓ��7=9����@���cF�qf,(��r����%{��!��-���a�H�^k6���ݺgg��Lo�XP>��DXb����[��Ҵ���?�*^-�Y�������|(��d
�� ����MD&qʯT|�2!�b2jA��ۭ��u����(��ԣ-ǀ�zqyM��f��$�9E�Z�� ��u���B�l5�(��a.�G��o���L^ӼL܎���䍭D�I�ԟ�!*6 ��M�S�*ٲ�}�lg�Qk���WZ�DY��+�iM�؁�4��(�]L�6,H�M�Z�v�ː��Ӭ'Z�9��R��9*H��76���~t���)<9�^�'1	�'3�PO�#��,W�$��QXt��c����M]	�J1#�^	Y��&~ dҰG�ě�Y;EH��Ӷu����/�2����'��Ԫ,��||@�nҘ=�h�!m,AտٵK�
r��I�~!y�u��O����)fVII��#�Y��[ K�V����.�P?��yq�Є02B�����G��]N��<-�	�cfY{yL!�.C:�΀�*�i��t~��Q1 ���I��߃^u�����q<��CO��S6��v�p�U?'3�_o�f 5$[�ӻ�6�>ᶱ�-��=�,�1n�ROm�����$juAh�����0�A�6̏m֍� �����,1�I
҉I�h����AN5��J<�v�>hDv,Y b��;�qЙ���$���} ����7K�C_�D�z�t'�xe/��y��Y(ŧ�_:�V�p��~s5~��)�ڱ�P���+�=�6�6+�;�9�18]��U�$G�%.P
(|B�(�Vr�'�ȶ��)Dr�j~aT�hU�#�hP^_?z�&��K<0��n�B �o�td�7;@	lF�G?&/�]\ A�F�\b<��o��y�M�9���<4Et�	zY�4�]��HӤ�M�.IԿ1�����e4*rO ��Rk�}J0)��s�ZY��sJ�`�����蓤fu������\Z�:�y���������<9�|3K��>9|����\z/s+����)�o~�"L<z*)N[�$����*�2��m�T5�����l�Jɍ��,��[�������5[��.���I�������1*��FsF\���9�<"�T1�	�`5K]�qQ���ac������U۩~�Go��� �S��!���go_��M�zG��k�����i���ۮ�M��@q��#pN�˺M��b�-\����n��㈂a��}_�!��3�Ii��8d���C�D��1�J&�F���LO��#Ђ>&O쿼i���Uhc�k��ʯ�ۗ�E��J���A]�S1*t#�����o��J�����)w��G�8^�>ǟsoR��~ew���c;,�\�A#�7sG�ǩ��"�� ��>��Mw�i������%שݲTu�e��iMP�7�D�sֱ�~�T:Ԫ�+s��HYH���
��#-�_�h%������6�JLb�@�=�������j��:(74q�H��%��ΐ�l}�Xyq�|Sjj`���YH��(Kd$�v��r~;�%gd�i��+��jY�Y��u��I��T����2��K�5�1������q#Q)��ij�`6��{+�Ao�cB �".N�$
{"*�^v��A$f�_�˼�r���P"��u�HS���I>�.-��1���f�8"+�&����d�N�!�:����{�T*�'��c�G�i�~}��t.�#���!,i��F�_HmL��[����OW!n���VI{��]Y��I}DԈʪ�6�J���BXjHl����me:Y�i�<�'�Q}p>��$�ţ�eq�wR�?��Go4�igp|(p��7[ �n�jѭ=Ai4`]�elVW�|�rEu�=��m%"_�LSW��_t��;�� ��ː��u�B�g�@$*MĻT>��uBJEȆ�M�Tr������h�L�{hC����=���F�蚜�g�1�3/��NV���T5��'B��f꿬���6O��Bˉq�u�)�x{:�
ԮC���fI��x
���̎��@�f_���/������jUH���>����O���;M�ǳ/motVn"
t��&2@F�W�Q!�G��ѓw[z(�U��؝}�r�k7���b'��a��l4*��Ã�k>f?����f??��KȡA���ʰ�m�J��n"�9x@��M���ov���k��Rs�w�7�=��	`|nҪ���K$v�
����_
gʂ���>9-��lp�m��z�֓�y\]��0T�yL��=6~�j���Vr����zHK?��a��b�@���'�&<T��%E���Ί��7
W��[2s�}vw !������tۏ����Ddѐ�uk].�G+h�B�wa��x���Qle�.�/���gCZc"��u��z��IH��)��@��(��ov
GNl�i��ޡ�0~ê���)<D����+DҠ��8f�n9=N�1:�$lɌ�s����ȸa���z�5���lUj�#t�����z�����$����ʈ��+��[�A�����ܦ�����V�'窈;FxN�%����ʇ����c�U�w�-I��#N#��b{�s�����є��G��Pz/���wn��9}��b�1/GZ�q$x�`ף�ȣ�����uS�l� �ׄ�!����27<��J���!�.�<F�$�_��X��`ws�#Uxj��o�յ�k�[�в��F#���zڹ\.l��8$~�CM�g윍�@����䠦�����x�ݻ�9��e�Y
�@� ��x*;o��#�i��ǋ�w)
݌�P�kk���8.��Ñ�z�,'q]���W�[,�NA��/d_��)�f!O���l�#���kݗ����Y̡��/o�;ȅ)���ؐY>_0�!<����i����KO��X��0�A�4����`���2�n0���ڬdŽ=��+���$�̯ �ϡ��P٧l|t¦(���`�lԄ5�BQ���M�L�B����ȏC!�Q�6^��fZ*/EG�;B��G���d&Vߎb�����5�8�oR	Y�K��4
l"0f��i�w�$��O��.��jquh%f��`b"�>�������� ��p�A���>9^ ��q���]����&%����ӏF���s�
�)s��\�i��ٷ�#���0N�T��/$��-/�b�rš ���n��i
��� ���0��\��^(�11;�֐���7�S�2wcf����-�1r.H��P���k����7x��j�%]���������s�^����6Nd�ޙgc���U�߸��k��nc�y`��?I#�����S~4�ǖ6�! ��%�%vVurU�M'XlxVHYEB    674c     5c0��T��xߕPJq-��R����$k��s���]��/��n·��FX��=��.���?�9.�9�j�qG��1j��6��H����eL^U�|}�F�P�ǮX��fJ�����~���y�a�zZ�����F�]]Z���K�ڽP(3��#-����/ ��#me[Ȣ�ofSl���\	���O8&�et�g9��t�S}]��h���n��qk/G�A���Ԛ�D���!��[Zc�|��rdO��������̫��Ft�@<�� �������nGΗ�8�qp/��^g�[��<K�ќ��z���y�1�3Z
[�^wP��B�#��E)1�	�0�BD>%��Y��8 ;B��O�"G`����#n����7�B���H�4c��6�X�IK�,q�1��2`�I2�F�L0-��I�!"��<d��:ur�tp.�_�97��]<e��GҘ�$"9�9�.��Ti��:�ZYNП0�j�&�Icn��H�m�r<��,�w������;Rg��1#Iј�7b6Ɍ=yV�Ţ]x�`�`
���Ӽx��_}�+�9FK*{����^N�'��B?�V^~X�� ���/X�x�-��yz�Y
�)}��ZX�S�Q��M?bL�Vs���R0����%|x"tG�Q�C	Q�<KkM�NJ�n��>���z`y��0{��gZ���p� lPp\�d��Q�ҕ2�}y媐y�n�q�V&k���p@�IS��x	�x}�/�6�[�O��%ǝ��	(�:T���t�R��<�^ZO��@FX������(-ꙷ�<��4h���?/�����{�����ܖL�_��G�?��l���zȤ�7�\+I&��Gg;$+�1! ���u�"QMYr�x�s���������ax<��|.��oi�F��gBH���ѯ���T���X�B@(R�Ѡ4�s��0C�*L]D�(�õ�[�����}���}��T*Q����FE��zEJ�fA��烗<p��7��%�C�7��z��(�	b?�QT��X�}̓RP0+��QM�P�i�������mS�9��F��7������ܧ
dX�-��a��18 pcd7�����>��\�Mt�7^VBW��\�,�>�V��<�u��Q�l��!"�S�(|U]_=���¾3�A	)~��w�A�� �;t����0y���ں$=������'�VP��d���^�v��U���Pg��$|2��&���!�@���SL���Liu�E�ViǄi��#�&�P�H�EZ����ASO�1�:��P|�!�)�3�o��l˴:�
#8z� ���
�-��H�1Wy{ Gcu��1 �s��[Ad�?}K�4W�_�Ȅ���Q.��^�����<�4�_�Q�#�5#͗rs��6��7��_Q��}I��vlc�b� ���+��m���ߠ����������,x<>�7\��0���z