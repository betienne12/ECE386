XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����!�?���ڢ=���)��;+�>�MF��42��o��C ��^�RmJ/�'Y�7���,��e3��ʶb���M�k�(]��D(�(�v�3�_K �]Cu��t�-M�B\�&��]"�$'E1>/C��M�� ��q�Ѡ���{�ET��W7�����vWV�U2�5$�u�����Z���Y�J�)Y'i�e(H�^5�)�NWǩ����0���i�_��r�4�����2� �r�z[��y�X�^����;�r�H�)M�p�6��o��K�9�x���Fe��A�l�i����5J5|�Rtg�Dǳ+�<$����0�#�4)�Ӹ
�G�ߠoј���.JW(1 �tH8i�l�8��ޕq����=zVWv���2�=K�N��@��r�5U矦LS�Չm���ߊe��H����,D��Ƶ!�*)yF*�{^,}qŧ"t
Yc+�w�,��8�զ�r�)� �+x��ɶU{����Ԕx��vI�7���ya� ���ͷ���]��2�JxA�K�^���t<*��r���[���,�࿫�9XF(!�¸�4�%v�	WL/��1�qz�x����:�&@8ʢP��>���i�6�q3Q�$���_C��#-���[G���Y�h���E� ���2�P���l��X��bx��a²�0��y��pM���_�ZM�Ý�Z�vQ�p����v���)���C�]5(�]!��X�Y���.YO%$ۂ��!�x6|62XlxVHYEB    9de1    1670_4�܄�Qrǵ���F���p���h���.��t�U��ٻ�5p�DC��b9�,Ƿ�׏s�'�g�Z��,��D9^�\� C�/���U�8��`�z�|h�? ����'�@������!;�*�~�"�;�9��+h!S0��`��*���@�Kο��<y������J�!�2��s�,�����X�C&D�I7�6|%y 1���q~y�GM5$ˋai���,�!��<n�P-C�J-�)@�.v|,���%��B��K`� ��
I
���m�&�h���8� ���C�^1fD`	}����P�{�6��w�@�T�nn;	�.n8��������P+���O��+XNQ�Mɢ:�G�sس��0�MW�0�{�"�.���&�����(d�ٝy/F؛#!�K�J��T����l(h��vs*+s\��I�>��g��-�8� �����O��j�	��v,A�-�P&�O-��\�ט����������r���i�R#ϖ�'��tb 06<5`M�>Z|bx<WA<��l�}D�B��O�j&�tD���H�Yֱ���>
����~s+�E[�U��7��.4l�T����{�QX�M�#Uy��hb���o��cg��,1��~T���L��gaY��Iצ����%�x)'��&�Up/�V�K��H@5X�D2J̲^ )���{/'��d��'����u� �5�9]�A6�U������e���z��S��O�F���ӷ�$�/\}��(��pH�Z���EɈ�k�&�dP�m����űڃ
]s0	 ��'~��J�k���JrO콉]NY�	GK������V����{�>���Yv�ٿ�!=�p��hC����n�bxmE�.�>�f�G}���T�
E�n,x�m������ΛA�����K�,Nzf	|C�QEZ�%��� \�`,�x���A��W� ��������m R`����c�S�톹��jF�ᗮ���Sv뉾0�y��9ٮ-��T�p���W4����h�A$�E|����#�|c�N���5A�H�������Ǳ�S��MS��攸`X'��U�����mH�e".(;� Nx�� 7?W�g���`��r_Ҁ-ֿ�4z̾�NǍ�[�)U;Mg�H��\J\�fAp�3z7OI+y@�(����0v��)�3��c��L�u@P�,�7V�zh�J����^7�݌Q��ٯ�~��;*h��I@yL��!��ƒ_!{c2���C[���lb1 �� �g��uf�c1�m-O�թ�v��о��P�����ޠi��4�(�?.V.f@j��N
(��VuKRFaM@��3���f�m7
E����H^�l��1^϶��k���S$��e�6;�җhثu�Z�\�Y��Gr:̩!l�J�����\1��>>�wP�3ۤ�Q2٥=uJ��ӍE�s&`+a��'l��d\����H%v��ɮ�
{Q�����Z��vÞ���L����&XjӠ���m�;��{��5�J`�F��#��tr�zY�HaZ��_����� �F�{�<�DZ�� IK�HhN�n4�q]�F!�^��l�7T�������'�ľ�/�1e���5܍�HLW���rX	E��/8*,����ʣ+QOP�	#`�
d�-\����Wh|�SlLd8�U������!�,V�~h6f��e�����\'�?�@�h����[��HܝU��3�jI�YIiF�ֆ3J�����嗚�h��ˬN��==5�����yi�y?כ3 <�E�rʐ�΅�Ra�If��b2�e��� |��9�\T11����D6�n~��e9���Mbym(P���>S�8��x6���/&�̬������:��=\��$Y? )�~2�vc���sY)�5
�<��2�8jR���s�ܙ�u��b�͠\�}�Q�r9#Q L�D9�B6��(��95~;��?2{�_T��_1���^@���(��rf�Y�L!n4�����TY{��U�U7����~�R,f�b�9��A1p�mZ2��R��՟p����"�+Bv##S:0Kh^�tQ�5�9@Y��-�E$chFl���xV���cS<�����ҝE�A3W���j9�a$�7����������f0Ɋ�p��Rq\qr��g�����(�)�*K0����*�%��͹�Dl����yu�������Z~OH�\���Y2�u����PG�jO:~[x �{�Y.��E�zĹ}���])�K�kQ�L��Q3m&�w*{��&>�B�܂�4;\UM-�|������sEv� �3�6�J{m7W�7���U9��^�h��G�+}��lg��؇,0�5��Pyk�HE%ڮ��G���r~���J���Y]��)�!u/��,�S����+�Mm�k�<������tF�l����̘M�Ej��W�m�|�كQ ���	DIN�.=���;gV��:Ր9�6b�h}M͌����A���E�fP��U��+\��Cf�^�	I��
����x4�ElW�A�{�
ҵ=�<�@�9�<ر�N�~�z�o�ҒK ɏ0(�HcWJ@?��:I���h���D��6�k�-��%���H�k��S�t)��a��pq��K:�꿣���x.��G�J��S|st�t�����҃���yۖ��2XP�$,��=�=z��嗮G��u�Qo�F|:�	��"2�t -���tS	5;Y�)��Y͙.E`��	��[8�x�ݝ.t���z��Uճ��{v>�2��	��ݳ;��v'o*Z��w��J:}5~=����O����W<R�r��ڌ����!�K�d-��_���\P߼di6���/�3=`�V�IB�� ��E��ջ��l��q��jK�˵\�6����>,̺ڞ�W�U��a��?$Qa[�Y����s�͝H�ꌹM�����H��ߨ�{ߵ߻Ua$j[�o��9��,��lv%d�F��w�)UVJ��v��w	�T~��F���V�x�IEɟ(���s����]��� Qx��X�����11�F�� �c�N�/�Z�Ge{;CC�[(p�
n�-�p8�6O;=e;c��c�W���:њ�=�y�h�}��!�k�����Qhs�F��Ec<��I��.����������Cԧ.�Y��q	}�n�D�ج�'|�����gX]a�=�j�$��c�*z�Z���Zӽ�O�e�?�+�}5����nH�ZejKC.��({.���k���4T7�}R�-�Z���ė
Xi�e�u�t�Ɨu�ť�1�DW��v���i2��{��h&��l.�;�� �[�<��XI�RU�Df�_�
RA��苕��!
���+�f�Kg�5<�A�E�U���1�`�S�Tզ�דH3�>xR�߻m S�M�7�s���<=��J������G�3�!�d2H�I!C�u(*��}�{U�-n'3:��	�{�b�A��O��p�.�EU��&I>��0�0�|;O ��n1:d��T<l����\�����B��UNm���3�XX�t�M��ؿ/���+fybݭ��{N��J��Sr�T�cAt��%`-y[�ȏ�&�b<��G8�c�L](�T��.8y�;Zd�fN��dUHS�eĐ) �P(/!�)�:�ׄR�����\��%�($g��\�N#b�!ݥl���R��Q�{D��q_��m �����k�l]vJdYӹ&S�,��&&|�d�ˀ��h��ׇ� �� C:GI���8�mFv��X��k�7�}�O,'L�arKUJu
������uX�R"*�_'�$л���-� ds��g�-��l����M���ߣ�g�a0Ж!~����[H="�H�(ۏ+sw�����Bh�ʻ�[�.n�n�?�6tB���W%�]�v������BuRv���2Ln�+
���8�Cy��5i$1O�v����R ��5����kꚭ����?�Թ�� s_���-�.��]�:魞\���K4��ę�;��~c�\9qhQy��
�1�j�ߑXa@	�6��<P�F퉄3�W���FPq�\�*�&�0?��V�z$B #o
h2+����[���Ph�}��{�"&eD�"6L�O�E��9���+m�4���1�a�G�	'U�ѵ���-����o��R{:�U�3�i������p��~���' D��̌%�ҥ�.����%�H,($�.J�T��)��(�Q ��e��10��Ixe�Q*�MC������F�5��)����?3�� ��/���qV����
��t�܄lO$� �V|�J��ؔ��O47�����q�c9(�k���\��$��_HW3E�_M�IP�h��EU�����+VJ��x�������ϱ��`�+(�A'�\/j�hi��CBw���q�1yUY�v󷡯�W"ڤ|��Kטm����w�T�v�V�c���V;�-Y%���э�Q� ː�����/�
A&���?�1�ҷh��`�����o����	N�G�̴5�34�̒z�*�k�!�T��0e��(��d+���N:�N��	��v/e;��.8i�'>*~`J��������'�{|��`�-�Q}��Xb#)�Ȍi��M��>�e���?�C��k�l�G���#}�P��7U�R®�\Lg�<U?�������͡e�$YlBA��KK�θ�t��6GH�\���0~j���y��{vI
��^�}uB��\71w��gy79<��z�]��/��Zcu�|�I"��=umM4������Fi$��2]��]�Ό�6L��=�ŧ|�Ѻ^�<(���^�� ��q���R���ٵv��ޝSZ����4/L���x��� �@�IWt�!Y4i*1��F܈�7�͘y�_k�Mr�0�B|�0�	#
�<@����(�$�Fzъ�8��������v��i�59�4�0�K�n&�۰�-��Ʊj(��#>�G�����C��J�w�^K��]gR�j�q��t(ge	&"��E<4�^}kPs���H�BZqSV�qY3ຫ���-377���ǣ�/yS�TBdp9��7�ޫ�-�U�~�(��e:5��^�'�	�`�%�_�����������m�4�z��uɴ<�r�bm�&�&A�ɏ�ݒ��9�ahq�K�'ﳹ��f�GbUV�ﰂ�jo��#6_s��U	۵/qd�k�h�)7s�/�A�Xi_a��`a���J�;^2H��Ϙ�6,�I<cyv:��'d3":��l��}3�RU5B[�?����kV>���W���|���E��6?l1xv����e^�Nk�k`P�y��TSy���B��㓳�E��p`��P,�/��D1�g���S���{h�f
��΢��
r		/�b�
6�UG��b�|-o+.*y��Ȫ)�����w=�^:�k�u�� -��`��Ϭ��7�VXj���Ɏ�9�k�d�u�f'unD�f��;zL�1�M�D2fXn���y�\h���~�QJ+�@_l1�C\��0J:H-���R5�_����P�O����̀�]�3�����F��+��%|�/�M���9;:�}v��LkݞvLj��o�K{��p3e�ڝ��]���SĨW�؊"�A��܎7�_8 ^"�l �����2�᚝���`q�U�����'�5��A����RC���HؐA_	