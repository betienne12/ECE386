XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7.��/���G�a��]��[-����]8�p�d 	c�&9Y�5�ٜ#Hd$�C�R 5D�$R��x\@�K�C�W(\`�
�,�Oh#��{�������mG,矮
Y(>�S-=`}:`�5���+�+��Ϸ jF|���3(8|Z	�����E��ƶ�ζ�v�}��S��!vF�tПYa� >����#�5�"Ml�'��69��|VD/�ȫX�;u�:|V�O�������l�Km��H5�j�8���%��f���R���x �aV]�zK��z:�ҵ���tI����=UB����sz@�])//�,��H�8���CaX���|����{-��l�қw�SD݆��M
"~�;�K�����Q����~�X�C\#.[\�%$�W�X�؂>����J؆+N��Q|v#�#gi�x�-���a�d;�J�K�r�\�PU����8񞔡�C7a)1z=��8��%0��c���,Ʉ5���[k}ړ��!� �K��*�*�IL��
˞Ǔ`�VVu-�������$j�\Ɲ��j�M���li��5'���ީr�;�X����6*�!yT�"�̝+2��c�mҊK�r� �lu��^����)��B�ffH����?��Sd�v�ز�Z�3����E�aS���u�^�:�v0-Q"K�][1R����&�z�VU�?���*�0�ݱ�T�G�Y}cj�q���Y֭���!�tvwpSd�[�e4��~��|it�}'��XlxVHYEB    fa00    25608��Fs�iI�,����2D������;ڶ�I����L ��(_t��M5�E�����@�S���8 �L���e=���)�f��z�89o�$��(���k&����qkR��:M���J|r�����0��M �U��Б�!���.�h��T����6��JY�������2[%��9��S��q ���g��K�m�I��}�� cZ�y3hq��(�A6��T��~�-��Y�rֳ.���l8����c^�͒n�f3:IF��ғ�p��gL �#8̹��Xb�u��@�m�+�7uM�3$��7����1�he7�$���5$l4��uH�۵�o_���cǾ�1���r�x0ԯ���ߧ��
X�7D���_<l���n��Lqj
H9��E�k��R�������5z�ݗ�*[��q�I̱��vUX�:���ԏ��Oԡ1E�bcO{$��X���ʌG=?�ۍ%w-\vf�o )k r�5�)���7J.��~�f+h�xA� � �Y��;�?���{Z|���Ǡ�����>�%d�Kڑ�=�y��D2ކ]�>����R��V��� ��m8�������Ȓ�"�F��)�QH�,��ϸ��~����tMI�S�z�#�#��y�;�B����RR�C4�8�S��zVT�6#��x��^��4$^�]�b����F?͛=�ga�&��s����<y$�X}�'��b�9�.m))�bq�51@[�y!ϖ�$+w���)T��E�<�Տ�`^V���.n�}8{�Y��qvn���o� ��r����#[r��e�`�����^�HB=O���G
_��J���Ȍ��}��m\�4�Ų��#H�4H�]�?�Yo'�X��'o�G��ne�d��uB܏��2=/ �(����F���{U@�}���`��yg�'��½bΚ�Ϗ�C�	�m���"_;�GNH��#�&�c��;��;���?�-r���o ���Ҍm��I��8�5��kjesRϙ��� {H��fk�X�b���G���T�@(���(;	����@7��{Qt��4�ҷ�OwB��[͐�4O+�{�q>��i�d30J��+<$�,i�*<!�������~&=����� !�^����S`6�794�ĩ
�B���7v���﫻ú�~�����\\��z�-�MΑ$T�S �?��ui4��Qi3���u��I��b[l_�}��ی����N�J�V���|Y�XY�:]<K��a�%�Z��g܈s�hrA�fu��M���;�%O�
_��:T9ݹ=@2��|�T�7�Q��<|Vf����Vzޥc�9���Z} ��G��| ���>����?�2��PO�����I���&�	dR{��dG�T^
x:O�������Z���󚺯$*MGY"弞�0:�_��K�{<��Z�T�'r������L�2�'�u���X�� t���d�k�N�qaM�!� �5��ō���]�~�!��Ǥh+��5��lt�ʷ����A�X�{�G�U�JN�����0�fcL��S�<�n����3'_��g���=��YCy�;�Iޡ>oL���l�	����C(2�MOyi����/hPtKo�~��̴��Y8�����{8��:��E?O8B v���t��C��]_X�y�ܒ�ľ����e��#��w�'�wݪ�:[j�����V1����UeHeu "�?��V8ū�xf����-+��e�cf�>c�,�QA�f��H��E#Qbӽ��O�h��})�
���y�e~���{P�cF;/ Q��$h:]�� st2��"E<ʲ��Æ��xw� ���:c!zJ,h�]�,8�W�K3|�%P�~{u%1W�z���opεQR5˕˞���G"�jMXQ�8�R�l;o�j&�ۺ���`��΂K�a�[?�Jz�IAD�4E~w�����4���7EG,w-��ǂȀ�L�h����:������]�����X6�B��Ƀ�0Ɉ���;�Ԯ��|�	2ƚ��4z��lɲ��T�F��+v��ls���/������Rr�fV����������J���zb�ހxמ�+����v5�~����%y.U�
ՖD�LT�@��ƺ�=��M�4_��}��sK�;mְڃߙ)Uc3�5-���_��Y���J�PH��A�������	(FbP�xOD���zT��� %��6�Rt��E���MN~�9,��A&��k�K�d+4VAݯ�^x�CC��E�?P�����{V;�dЋt�̂�rN�M����03�,�ѷ�g�ߒ췐;~���]u��Z�z�>?��ƽ�П�Ol}^��467!��S����N���=%K�V�"�a���ʎ����r�@�lS��|��v- ���$67�����K7⽶W�i����Z����P�ޱ�8.!��"�*�(�|*�O��G��/ŀv�KA�T��U�BŁ^Ɖ8_ .]b�7<W�'-�%8ᅤ�0�)��S핻>�8��|vh�&��4�_� �\��z,P��@��R�$W�J��~�ƾ��Ħ����JQ�B���I�o�<�"a��+x��^�v�@�k�Î��ӡ�ɳ�+�Lu��K�px*���n�2����]��"��Z�li��e�!e:���;!ӇI�&��+ ��r���Z`��]�M�<
`�U
d;W�HĴ��#ۋ�#e�Pi�r��	�
-�_Ub�,���]C�l�uf5`v��]ݍ�.�Wѹ�ׄ+~d3�R���o�%[�N���bmc���GPh��m�(��ݵvQ�t�8fz�?6O����y}�6�{x���|����g��V)�	֐���@$^z�3ﰮ��RZi	�~-��j�^���,v�-GI��Q�����$���"�x�~r9I��$(�����1�Hs������_��Tp�N�"�m�� lʐ�\c0�mT����x:��6[� �e�N��Q�(� q���Z[>�G�G��۰���g��J%Tn��/��P���Z�b-��C86�1R�94��J�>��L\�����h捍���>6Hj�x_lTO��}��?�����J���.��=����I������׽��h������^�qD��<�0�%��WR��?dC��]�}�|q�߻n>A�"�U܁�S��Lp��ee�LYc��ttF9(G�̯a��B�����0=�Б%F�m%�|E�h8�U(m�� ���E],+eh��D�ɍ��.���E~�\f�0�4��"�xg���̟~��
����ܨ$X;�B�V���V�<u�t�<�N���-~9`[q��+E�)m�ӧ"�*b�#>�G ����D�(��}�:��^AتԆ-�d��5��u�:Jy�@b���T�N�ór01)�I�V`w:56����$q�4�3�l��2hf�Y�,�|�����r̀��&��k$r�O�� �k�P����3j�~zqn�=C'ó絵��0+�֊5��1^�)��������S�LV��k�Z�s�4܍?m�����9�Y�Q���;�$w�z���?E,�Ǯ���;�sZb��S��(�D ���/�U���4��ӻ'vR�	�a'�4�>����ael�w��_�ҿ�AM��͕�K���|�S/YV�fL(8?�QV�!A���
���G+Zr^���ʵ+/L�t��8�O���u�ʵ�dI-�:�n�@�&lջ�J�v�@Œ���+)�� �ע�p���q
E&`��Ϊ]H��:���U+A��l��1��� d��K-���&K9��l��,�f��"R�\��a��T�c?�$y����w�y&eh�5V��s	�~	i��@��94�$ ϢX�^Gy2ā��5V5^6��:D��l��{a6��ΰ8���m}| �����.�&(s k�z���/�-}=W�'��+��'L�ס礂�y�%33D�>8����6
�!�
��L��L�"����:�d�)�J� RT�6[[����Z,�I�l ��}7�~��Q��ǹ>/ �,�b�&FP��س�<Ȼ5���8�^��f̢L���7ã1�p�����з�ɜ�mT8���v^�4eR:���$����'���v�8T���'��p�º�,u�gi�����I"�A�b�e���������X��=�m}���˪��w/U����N�Zv�;�����:�D����jiUp �IxGe��W�C'<��/̭�l0�R����Q̰B8H����΃�θ�5��NHǩ���j5H�t�m�He�6�̚m'3�Ȭ�`!4����u0&�t59՚H���v��<�$3"C�Y0a&�T�kX���Y#�O��nkϝ�ۀY6�	��ŬY���&J$�W�^���XF�K/�=�����Z�+�$��a�.F�Y�"Vb3������>qP"X�)[?�C(�\�s�������v*p�I�v��>����
�(�wb.ݔ����R$��W`5v�q���U��ɰO��TVp��ٟ��RU��9`g1��T�,�r����V�6y��ș�܆��P'Q*/�f�,a��� ��~u�^3����K1��fI�"~D�Ht������FJC��NM܋$�����&T�n˖��=���.��2���A��}|o�=���.�6����9.�R�����ؤ����C��cP�,����l��`W�`&��I�=��w_����V�RS��J�'����e��{��E8^�W�̪�Rv��x�c�ŵ��Lj7h�]j�{�
~:!Eq��q��>m�Y���lC#���C�
7���F���z�a���Z~�MThq�(!���a;�i2;��8h�bf�j.=�Yv��^�M��*�ό�Φ!m|2z��m��W������B��#�Q�q[�YZ^&,s>�<T�����G-gB���~$�/A��FKrb���<���0�K�E^�2��NT��VL��#ʢ4�~ <f�t�sפ������\�9���x�x�L�Ϧ��g�4����!%���aqJ?n@��K�U%�++��NJ��A�LO-Ov���lke��cƠo�%�@�x󧑾�Z8P��vLE�#�\��38�?ô��^e:�Z���Bڐ�D���"����4x������R��1hQ�<���!loܚoC[�A8�x����N�C���j6�Z 4���4��y�HB��{m�[�xml�_�� u���^�Z�9��X�a ��P��?~� F�$'{K�!:�Z��:g%c��1�g��Jd�e�tֿ ��-Fq�"��+Lf�*t�
�A���>��8��&G�ኴ��Ix�~�4~)�x%Ĉ���ݠ��O�!祋ע�ߵT��>����6h1x����sH �>��A�V��Bo�4�'\������CC��^���?����,9�|�w�j ���B���:�aH�ABC�"�*�x0]�_��,߲9o��G���VN&fSpKm�C���R/G6��,k���z��Ţ���n�/a�XR��|>:��6�,�~���|f�̹HP�ˎ�F��܅(<p��H�D�6��m¸��q�;h�3z$YCՙ���܂����� N9lS�W��6� r)F-\N_��X���gxv9�y}~t�+ҒD2.��(z>��\���� 4,�����r�wZ(��53�ҙ�q,�a�J,��.K�d`�ũ�(W���ڼ�J��^᎜[;e�6�����Jm��Y׺I�%���6����	�٘��+�7�ڈ�=B.@��x�-e�ɶ/0���*o�.Zt׹�S��l;Y�\ݍ�cӏ۫l������,`g�L��E���Pt�E\�Jl5-tf8�#�1�Wo�%M�j��65T��ĩ̞:M3B@� ��R7�$�i0g����>6���D��rҙ�ft7�gjJn���t'�b4�-��\��f+�="l ��Fh'�F���H�n.,6������cr�W�A�~&�-)1[*�x3�V3�Y�aN���;z+�	-/���|Lbnmȣ��3}����cqy*����T��m>�آa7��R��؄�DBc$�;u��zV>�a���R���0�iy0L��>����O?#h �a�>�+����qZ���
ܔX5%ȥ�)�v��\2L<i��f0�c�T���<��BꇐN�z���-��%�V�<Md.�̩��F����~wO�г��ٲ'��-��g�������[nK�����f��Hw7���6�s�FL�OJ�É�^�eG��Æ}�r�g�{\(�7g����d4�؛:۫~${?̂�$���PEv�y�v.�4ޱ���d?��L>sʠ��Ƅ�e�#[���S�6���ty<���.�}W��]���N����((��dL_��gv�!��^`��I 9�G��:��/����J�y���6[�Eg�=KK!�A�j�yI������	�}����6;^#͞��jW�ꓫ��g^���~uc���R�l,慊��Ÿ��i]���[�豜9Մ�ܸ�45`��q�I����b�ظ�iFe2�ia��} >7��t�z���U�L1�P��z��'(}�x�3^I+B�����{^O�?��&9�K;@���i�j�����	y8��P�*ɓehbF��^��$����T\����T?|�H�%����	[��vI��Ήf˴���x/���&M�iĶȶ�?�}Þo�Q!<����\ͫ��A��X:"��P<K	=���gG�-�9naS�9��
��~�/�����pl��h�#T��*�4���~2OTo~x;�d����_�0^�~	|�	�o�B�_��N�p��S�;Ov��ԣF
�F���.�<����I����9@���¡������a�(���B�$���N]N𾖭�e�gI�V��B�W��E��6����j��#�3�y�!�6J�/�-��2�<X������u�d�,3u�iVQ�V̩�C,Խ?�����*h/�ܣd����R�Z3���#@��<<JI.1H��eL0�e�a8���#99;=���Bo	�7\T���ֿ����$�Y R�Vo�8�H*9t*�J��SY�)�a�yM=S��A���F�	c�N��/�?vC_9�I`�qѿ�r�� �GZ�i�v֢3�J�n�s�"Ԫ��]��i�G�[4�}�jMW�\w��Tb�s#��LA�!7tY�4�iUᖤv�����;v�q���7U��������/��*����Sy�v~�v3=P<wl��۸��q�U��;��i���ɋ������p��FP�Ѐ�vT�fЪ6�����i�`����s:ˁ��C3����۰�GE��30U�)�z
�i�L�ݏ�%���h��Q�3�)_̠�������������:�Q���/����v��|R>q�+ &�����CiT�#Yǻ]�k@�؈\V������u�t�距��3��D	c�8b���k"���#�[?�M`��7H�]���Gng�Y�Į�
�͚�ɫ��������s��ve&X�Q�@�vҖ��$,%u�;�>M	Tf�h����{2Vd�l �L�V�N�~�`�V�4G��oğ���ylwQ"n����w�%#�-.z���1�֦�Ɗ�-}eP1S���jK5�a�>W��m���		�F*�&�y*Hu�}6)q�Ɗ���X��nyJp2̀��i4Y��0	�h����4v� � ΂-�3V[`�x���+���/)xc{����i���lowp��]�����i���E�G�QV�<*�\%��f����c]�1|������$��&<�@^M�]�T�7�$ǿ�a�xL"���Q�m#39�8HP�[�*�!�Y6e��%�)�������fL+���p�V�v["��\��( y��+xr39Fԕw:=(|���Z�qX~��z=�.q�uk��J��7*|-�MsQ�6�j�F.��\�{�[��U�� H�u�U�!���\�%��,�A����
�GxV2���s�h��5�����J!$�����Ă��Ê���������U�@O~��<����`�*�4(j
�S�(A5� ��Un��,1fy����ޗ�G[��f��x����ej��:nR��_O�G��P��a=�g;����0�l��9z0(9Dl#�4��K��F�g�eF�xը;����AoѢOɐ2]H�a*SoH��f�uG�V������5�?ƀ�Q�Ny�4�0�x�%�:��C����d �>�_=Dg��T���wݾ�Ѱ���/~Aϳ9K��e�/o�n��I����$?N���{k^ᥘB5��d(����+�\=�´1���(Ԭ�i&�Q���+�̮�y�E|�$����(F�=F곎�c�i�iMpGC<�t���=�g�.b�*��e�s���zB��h�h�	����mN��F�I�G�����-�֩�,�cyD�VeՇx{E�l�ZU�~��W{�����«�^H��u�uv��Y[ј��SO�7�ᮺݎ����B�l��K�ӌr���Ƒ�]�e=7dJ%ֶ��֊�o�:ā��'��U����[㌐�d�Ro�w�+�!Xr!���t�ʇ}�%��A�Z��O�!�$w��щ+�MA���iY
�����e��ف��i�b�lEF7�ӄ��'�� }#�^�O�r�,і>���~B,��>�Ф&-�ig2L�ܟqS%cY��]���Ӑ�c5�գ������,��~�`��>t2Z����:Iv�7 �۹ڻ}<c��9PK���)�@�������F��"A��Z�Ӂ��_2��:����i@�]#�ڎB�H�3�f��NC۴�U�w�M/@�K#��GD2ev�q�^�݌�2�����6�OaK�^�9N��f+��O�Kj��B-�t3q���ZE��$Y��m�YW'�Zu��-�}ƹ���T��$��=�?M0-�ak��&|G��]��c���R�5�ùè���.���^�wi��xGߚ�^ڜ��a>���h��%�L�֪�L������W�ب=�s�
���S�"���;,R��9J YT7:9�A6��������3Ⴭ�=*��j�$-[M�l �Dy�k�AS�	�nu'��rxܩ�Z��V���K�Q2:+��q���-��!�*h�.?&�G��!~��!�r��gQ�g밾m��ؽ�!3��d�+=?�*ET�����'|"M�5 |�r��/H=.��l�+M>ܣ�-��K`��o5��͂@L�kgX��)H@��7���\���{㟰98� 8z1�	����i� [���M��*�r�;�6��v�x?y�����=�MϬL�ٞ�J�Q�H�2|����/˔.�ʹ�}ȊRR�pSmssv:N��8�3�<MJ��Fh��U��9^N�{_D�v����2LE��#�kS�c�PUk��3� }쮰����+Tp:?���t��t�[���XlxVHYEB    fa00    14b0u �g�9�������B����Ǹz��Z�2EQO���|�.��ej�U֊Kb.-�Ut�4]�<COVK�쀘LaNc��g��ʀB�+o��!iu�fHK?w'���Bl^�9�.Ӆ{?o�|�x�r��F�]�hM3��ԛ��\_�e�O�a-�"�W��H9�F��0SX#L��(�X�M��Q�Ċ%Ǿ+����߈L_Åݾ���*E(�w��H5TY7���EOz� Ceeh����������_��Xv���h-�?-���xc�X/%ֻ[����	%B�p���S���d�R��`����U���+|�,NYI����n�}�'FN͝1vS<yݸ Y~aH��u�Y�bK,3�1�M��|�G1aEq�b����J٭�K=8�b z�߻D�7:B�!
N���tk��:D֍��r·��,03����-��'�SF6y*G���"r�Sޒ�6ູu�B�,�x[�|�(D$	��t@�1��. ���I.�vb�(Z���u�k����(�g�����b���`����|���Ytg"as�`�l��@�1h켢5�r�c��fd�����y~/K�����P0���H3��v���2rې]�����\�q�#��T_���"��2JG�	U���o���*����P0$�0I���L1%G7s�7ڼ��3L̢�'�O�)HX>Q��jJ������0����{�D�!��e�buDY��ݫK~k֦|A��ݓ���}���QTc1j�6�1S�@B+M�U䭣Ɂ	W�/��@Jl��e��Y:���R�4Dr�C�� ����j��/��Ғ�R�3Ҫe*��=ZW���L��:�����=����{Ӓ�j���VM��d�D�o�{�	��=4h�uSX��ooA��( ���x`*� |��^��N����A����,%Ĳ>5/�/?uy�BzF	_ݪ�u��ɌEC�z5�a�:�l�h�O0n�WH���x=)�-ԩ�	��7?e~�R
,��ߢ{P���-X[�5�+�]�����:3����D�P�p�ʾGZ��j��?���&�X2&��=�%���ىqȼ�2�7�&n{�Ζ$\P\�Tp͐����+�	-@����H������{������ 6���%]!�(12��;�R.�Uۖ�}�,1��h�g�ЫO>nD�y�����d�Aǫ��dxY�p�>�>�(a��S�Ibr�D�8���e�{J�i�fQ��e`a[!Z��	�]Z��n=\���o�!W\Y������)��ӵ��.Ň<�Q���0��%Ɠ�溚��9�W��[&�ş�s雬<6H@��^A��������m+��� ���Af�'�4j�ǃ�WS�Ƌ���ytt.v����;��š-�nR�v�*0���x1���� �P��wf�&ٗJ'T��OJ��-���+�{�b�O�mI"t��J~ţ�ɇ���X" Թ�Q'�?�����8]rC�n40^���N�C� ��o�O ���V8��Ne <kD��Wo�==Ug�'�&;gع�j�u*��G=?�ܼ��ܩ�h�y�|�2�u%9�|mK}5��n���V0IB-4�ۣmg�fヱ\i}"�J7 ���1J��Ȍ
mށ��pf9QKN�H~� �X�Ɨ>���i�����C���\c�ܥ�@@)^.�(���3!z�K�J��CI���@m���'��竜\șY��г��ft�
�����It�7��<�6���O�|CXi c�à� y���(]�1�"��8<s��;6/KSƈ�Z�"*l�Sd�[��NA�g�ν�ڤ;,%����]S�\ a����~P@j�;��6��Fe1T�}^*�JA��]�����V7�Y�-�N]/���/ٰa���f(l�����a{�!��׽�}k�E�4��c�saN`OZ����ƅli���/�W��L�Y�Z��2�y8��wa{-�8��N����K�	{������<E��$�� �������>�h=�s��hU�.Ǫ�0w�s2D+��1K#��B=9�o\���L���+��pLn�$���ʡ�~;o�q����BY�5���L�xə.̦�+��������u�Cξ��@��{�c)�`3@R��+&2t�+'����������[�����S�F�ܜ�W�ħX[����c�.ʅf��7��x(a/��m<_�!�v�a�X�F{EQ��.�:%�0?T���p��t�t�{����/���8���х�<(�og�Hu��SF�N�d�j��Zw;�m�r���T.7��e��7�P����u/���� )�?��ͦamN�]����:Ԭ�ȉ����,�{�H9+t�����R����Dݵ.�Ċoۙ�U�ۈ~�`	����;��X�]Զ�͌���x�}���i�Xj`lMT�v���F����� .Kl�)S�0+Kލ����G(|���$��sV�>�O��m�l �(-�������S$�� 3g�$_ӡ����[Р�S4�]x�`��s��Qh$�:qA�_Y_\E���2_����A8xRp��ֈO@`��Ԁ���Zi��nOJ}d0xgt�ph*'-I�ݣ��;�΍lYl�"�{��vH��ķ�&��1���]X�Š��ҙ�Sm
�W�q�jP���ؚeD����.���{b��ގV�h���.�<l/�#B+�k~�+ϭ���V��tP� ���F�3�9�
^ ����GymT�v�nB���&p�4,W��Cd�`DM��/% wϨ�U���D�/�ҳ�"�������9,�ݿ9�����A��.�5k)�V+���^�9���ϑ Xc�Mp��<�+kׄ��A\���b�`�@��#�5*5.q�R��^��ۅ�}{L�L�{���M'
��j��s��H��n7����]��ki;�\pe�4�>�p�]��aC��Dӎ��x�8��z �)ԚԢ=E3#�3{�9�+OX��.36�W<��>k^��/���}	<���:������� +y��@如��u�GP�3�[�>o�K.'N�/|������o{��%�	�ە/d~���3�zjy:�; �s/�W��1O��@�<P�X�+����n[om&5�L~m�Z����"m[���_��.�2Ҥ�B��)����~ E�:V՝�5��<O��E�)_M��sЗUwF](cB�� �aj�E�f�_�A�N)�"���1	lV(O���{�/�eZ�0�����5��n[����r�X(��<=;W�t�TQgt��T��W䰇�Uk8f�fЃ���� ���k��#3��9���)�V�c$�S�8��4�1Y�p�
��N&:���(!(�Ks�Mg�&�:_h�'s�q���倅����Aj	�� ��:*2.�-�+{� ,U� �Y�9��[��#N��R��SY����y����f��T�K>�p��Y/L�y,�<�)U;���iiG�����C�gg�&�UZ)���� r�F����#2���a��=�q���� ���Vnu���*B��\3`���K���@���۔��tMbVY��4R�:5���="���w8"oYE/��[M�*Cw�J4�X�>�
6�0�j���_k��4c�݆4q�ӓi� �?��	����V��?]�e����ЋS5��5����=a�O�G��1r���[��0EC��J�`,.x�Z�m��!����܀���/�	~��Q����Cg=?������D�@�#���ɻ�t���7�2�j}�<�(۶�
�����,�A�0���/c�����8M��~P�)u
!�id�d��w!xʍ�^�YS�m��<�&L�%]��Hq��x��A�3�4ŗ�?�n�ی�w���I�������ج��Yc~M[�t����\���ѐ=Hw�"�?ǹ=9G;%�"Z�8��TŌ\G)L~���g徺N��xQ�}�!%����	W�Qm�3���L:į��\�֒	��u��ɲ��d���	�9b~�p�����9C��^�%��s�3�h��O��G�qU��ˆ��&��4_N��Bo�|����e��k�U���d�/���%ڠ�Ͼs�o$��mC���a��K=���)���1�;M=�\�:��A��$�1L-]�M8k�ȿ;���.�����(����0��j5�|H�����W��d~��M=��L��:}h��B��Ҭ@U��_�%��ݺ:e�	e�u�g{<�h~�_��
R�aY�Lu�E�ϠH8iK"Ɂ�p	L��]��ƅ�6��\�a�I�Q+��}N�e˾Ek���=�̆��'l���-6�̉3q���	��$:W�bQ�m����*݆!�ou��J���c�~��/?J���S��L`��:J0���'��ǖ�\	�M$f^:l��r�E h���N���6�s��|�P��pN�M�&�a����Oؾ�n�HY��dI�7�s:���G#%+�������yp�l[�J�/�y[`:���-f�T���_QC�^x�"m��vkƐ���d���d�0��0���D�r�$��� <*���h�o��;����1z�}�ϋз��$g�Cr`�����hC��2��H�R��4P�.���'T'���>���&	qPcj^t�9�D]�Q����c���N$Е��u9�4��]��{�\�Uʊ����MR[Y���a7�zi`G���b q�Gg�jp�Gd�/S<Y�87���P����L[�#����m�&���6��倳��_2g3��S�om�gՆ�|<3�� *{HW<��m#��V���ğ�xs�6��9n;�Tu�Zg��x�E`����j�>�L`�A�أ/����Ң��1��}�hS�r��[������h��c�	�,%9��5��	�nk��B�%?[~7����&stA�R8.ݷ	�#�r��.H�Q����h��X1���(�\ꩂ��V��Խ����7��^������Z�Ȟ����/�a��<&��?e��t���
�1r"7\$�������F�],���we����P$ &�@�`1�xx��$��7��ݞ#�]ϾN��Rdu�pw�1vr�D���Asm*YAƥ�����j�-��E���$�5	XH��a�6�J�4�7�쉾�S|V��Z*P�l�29�i٦���۱ Kƛ�i��D��@��>� i�£b��c�<�XlxVHYEB    fa00    1880�� �����X��a�1��U3ʊ�M�n=��68p�YؠI'5�|�!Z<Ӥ�_����{��^�<�S��XD��w����ƳM�
��b@&;�9�b��:�o�ĤV��j±&�eS�׀4�L����..��n��ɒ@����X���
�h�0[�z�`����44+�)�l��sվПRө�~G�0O�6��T]�&�l&�0����e�[M&a��M��1]� s�ǎ�������D�QW��"ց4-!��d��[9�P��������\	6B�`,�_4;͙�{�L(�W��O]gz�+D�g��kM��.�t�B㛰���"�U�-A�~���X�����lK��c���ϩ6^`�FM����x��}O7�$�L��Br��2~�;�e��"��Y��3
�]������9=-�ݚ�p2�_�.X�q��`K���j��Ҷ�����)������<Ҷ�S��6r�����#%gw�{{��a��p:���=+3�I���T����e���gg|k�p�zB��,�1�K���I����A���q���W�Θ3�� (,Ӄ�\�������Ke����k�R�MY�~�N�І.�����Y��Ě�
�5�.�m�7�KI@bIF-P����
���P�q�o�)U�;j:�!�ZpR��-������r���(V�� ��@W�]i~e�C	�WqH�4\�dϑq�%����۸�wU�Q2���J�^�����P�V�
���@bJܙ&j���jW�_�o�GG�6��iڶ)�1Y6(T��\xЧ��v����{�R*�tc�r��?k�����vp�jv���le)���L�-�I��?����M��*���wZ�3�E?�ש�4�n>3u"�#��\�I~��H2K�Xߜ�vG܇�Er ��;@o���j=�Ԋ^��c��p^�g0���&B�w�ݥ��h@5��tjY,��	�2kR�5�b�r�J��vHS��y�n��𳝘�9��$�� ���v�32a�O.8I�s���|�b��o��[!K�81O��|np�i�il`��9P���6��x��q~�Mo�4q!��"�ꋓJOA?���p| Ȅ���E�w;��iS��b���y����*	��)���cy�Q��@��� ��X�M\�_e�#�����v�ƂS�@����y�8.���S���I��R�a�)���ղH�yk\�`��:��2�C��ؠ�0�8'���O:�ZƵ�MF��	�	xBkh%�Ӥv�*�1b�����s��-'�j�]4��MV4��`�B;3?o�$�:8M[ٵ\.��F����o��xT�o1�r0u>�����ҥ����ަ�lY���:���k:�ؿ�L`y�Rкp�TY�H���8�g�i��M�?c�&%�� ��Vb4C4l䌤��?�Au4Qr�*�r}@'Ȝ:���e:
'�G��^�{b�en��C�cvo��U������v�L%o7��ƫ1܌OSz��0�n��"��v�~#0��S�G����ev#��n}9�q�tH�V�s@�Tw�g����>!�Է����$�w�X�tb�2�D�G��	�o�#:���~;�t��|�i���5KfŪ	��ґ�ek�,$:��ǜִ8M���d���;y��J<V�?�x�F��6�z��D�V�4D�)D�J�hD�La�L�C��Ѥ~��VO��H��UO�5#f�5 W�=NZ�;�/ܶ������p�ѳ-Q8xw�X��۫,��[���	�����={��UV^��C�;�feť���Vl�?mJ	vxd?���.��/ΆN�hDE�4���I�8��n�)b�+W�GiHǯi%	��5��5ܧ�ӓ]�C'{��PN�⸡-4�s,4�-E&׮���n��$ԧ��k�Y��k|�
�)��BH��n�ڮ�{b�լLͭ��!2��z6��hA�WTtE^���<�T�v��K"����ﲷ��{�Q��J<kC�ڑ0���@��[
N�aq�	�B�J�u�����S���]��� V޴4�"`3UXjS�����>J��.�r.c�H�W����j��̿�;�0�ĥ�tG�z�k{_t�j7����e��������S�)�{�Q��t�S�$� 
%�e&9�l�d~������+o�.u:�B�H��$�e)�����!Z��%��;���[�����Ɣ�Q�Ո+�hw��3K��T�?�E��<��y�n�[�����p�~���\�t}��$�C�:���>�>_�~JţJ����N���7S8\6���g0��hf��v������<[�`G,h'X��m����53"��Y�`yPz(lAP�����\Ҫu�SCO��������+�:b��c���� F_a}��
�� 	К
���*�L�%m{�#2S���g�ex�TN$�(}�B��x"g9ta.y�J&�HJ����R�R,9��ؑ��>F�)�g�����J��#G��7�Ӌ��r�YE;�v����L_b��p�-�?<鋎%Oz����(D�P��q�;�|[����`�m�l�5�YT#D�����e<7��Rx�0��}������쿾��\���Ϙfp���,��9K�Ԭ���]R��� 2��=ς�J��������l��N	��@��5A U-��y��7���^�X�h�Şii���]z����V%{�#��r��+�r�1��$�A����J���X�.�Ǣ58�ر��U�A#���A�H�]��k~�=?�����T�҇6��t��y5��&r��E����}���kܳڋ���f�<��b�G����A��-�ut�� �2J��ٿw���9����TZ���CˬvJ���<* Yg�m@���K���#�US.�6��M[1�;3y!.C��Ô�_j����%9��j)��d%��ң��P��f,�~v�qSfV�C<hO�I�2��W/"H!�xQt	b��	[���M��h��&�m��m��C����bn���v���_С@-Ķ�_�Պ�T��g-MQ2Պ9��%VC٢�+���u +*mb�o�k�?\��\�v�)�6W/$�)I���:��95���� v�<�wS��`��I�]��K�s����Z��(�+�|5�;b�EF~.n���fF.3�f�cd�$���
�7�����$. ���۲F9=q�L�8sR��4�(��1���	���{��Ceľ�HkE� ~���	Ʃ��5�{
�;](0��G.G?؞K6���7�;L�9&$�K�H�II ��?b6�W�5M�0b��6>i�r:�r�P%$��B�̮�i�J\�����pXr���X�o��f�f�}z�4���Z��Rb���F����dVSz�}3+p������X����?9�j��Ru�Ī�JG�6e�/#��6_\R3� ~�?���I�^��ϓ�&�g����f�_��+鍍� K"/MZ��@J�hi�Yb��`�r� ���/Er��^���߿�U��J|�PXH�Ը+�i�О�-��w2�<s.(�u'�W��-�eW�͞�[��gkȏ���<8x���I��H�1Ik���¯',�h�-#�����z����Źc�D�%��.\5���}�$u���F�z����X�[�) p�Ŏ/('
��D{|�&��Ȼ���T�&���d�4������8��+ᢵ��U	�B���3��(X'���%5t��|��S���G�og��	q=4�*S�j�k<_(�.��
+e�i�� f��\�7�P�����S��t����w:���}�����	�5�{�C�`/?@�|S�>��!p�������#��e�J3�̆�RO�����~ �z�����w)�ܿR�J�̻o,Z�d����t�F����,z���R1a~�F�^�'�F
�eF��(~��F�/ ��c�ܾ��%� k_M�O\�P~0O��BҞ��O� ���2v�@m�I�pq�x���Vy���J*�v:	|�����Y:�N�dF*V��8�a�Kt�6Id�3���^���V�L}�ǰ��LN���׽�t*��,J<*���|a��J�B�@tč�r�X�5:T�)m޹�̬�'Фv@�[N�&�˳bp�E7�N��*��I
N�,���d��=�L=8�ܐ��DR��Ř)��W����6���V�@C���,Y�`��@�9z�]��in�#��D��Ϊ���k������1Y�-�+A��8W�c�H���y�k
Cւ�x��˿8R;��g
oH������}�;���*z)�����:�xwR�q6���H�u�*��m-iy��9�eS�`�q�Ϻ�8Ӆ�cN](j}=EM����z \��A,�r*�/����RM�;"|�[��v�}�>W^.-ǵ�N��!�a��a,�O��h\��|�������v,	>W�S
�w�3����ڑу�IP#���d�/-O��dT���~�?��~?2*c5�H���*� w����3��>�[�o�w��%L*{g��t�\P�d;}��������4�GD?�>Z���oqɣP��Z��Ƒ=F�������C���N�`zOp��S�҂�: i��U�V �_��,�/D��'���w�3!cJC��o���
v���eu��_�`'�[e�G�Ri����g1�El�*��(X6ѓ�:�-Ar^4}��q.iF����S^as�6���M�@ʒ�D���+� �z2_;�	i�;?��#S�O���c �&Z}�tG�f��Z�����i��{Yuv��`�	�_�+��OuROkT�>�MAt�6{̹ l;:�����\I�Y���iA��u�L�1%mi;� ���ì��7
QS����J|�ɡ��((�N�;p��Z�8_�]k��7��?|�R�n����`��ƭ��Z���*f�B>�QP�m�~�1*����� '~s��qM�H@�A�߮�-�H��^��t�C���}��G��Zߤ�^A:#Q��ؘ,�ᢻZǌ���V�R�(�w�� L�!����F�t9���<����i����v�8�	(�������0�w��ǦX���<_���RrN+����3�0�4�O���یĦ?2$�>(���a��sC��_��8G�Px�U4�9��"��OM*1���|5U=
�T�c�0��f�O����owP�@�	��ݏ���iCb �T�����x!I���΃��N�@7�F줘I�	k���`�����n�ء4x���*��=�4���~��T��6�f�S(�U`=mgl��� jo^���g�+*ε=L��<s@��'�yV��ȼk�+����l�d�`f���mY	������V4K�Dp�%��m��.A��OĎ��H���T�|�6�Z�T��w�c	ᚙ��z�%�ӍN�����������&=�J��w�HU���%~Y:�ǅ�:�X�#�o��Zk�k�RZ�l��䖨&�q��JD.;�:���W���b�|�&���Zj̝��"|��QK�b������d��B�e��urK�l�]� �"��;�0J���޺��34UQ:B˛0��m���a��B���ͅ�qb�a��(a�k߾�ˮ�<�IR�k/t߸>2LY�!�6���Scx����9bQ�/v��\L��R$ݱ���)j��	�\W�S�ЂQ�	}T`��8�=L�@:�/�f�V�����1F7�kƤ��]�J´V=pY�G�;q�t����S߫����k�(��'�>�;�=�gt�v���pS>�ZO�p�5	Vʭem��_ %��QW�'Nzl�ы{(�^�����:�dc%i(�lͼh|Q�o��+$�-�K�e�[b=�؇��&�8�9�u�>�r�9��+�X�;l�p}(��Fֿ���S���s^�B�q���6M�#h���n�>%��}^���hGhY'�e]7�RPm��ݽJ��?Q�
���'�^6;�̴�Q�X���r����q�C͓*^l,�b�Q�5�^+O�o<P�{�{e��t~��Mqv�l\n�K�nT��Y��p�8Qǉ6�Y5��S��^��C;�WX��E�ФB�z�h7���;�  {=:�,�@m"$��+������ִ��a�3w oRQ���'�]��ҿ�#���t�b��7�Jm�"�y�EC�fXlxVHYEB    fa00    1910UM�Xր���Xw��h�0�B���<�K��������{�̦р���R y�f���?F����b �瓧�a������^�~����l��pv���V�ϗ�Ə�W�_�� �OR
��<���"�6�rA QzN�.��ɤN���Z�2��]�/�[�H+�X�dг�8�Ţ�	��7�crx��N�-5�L�mv�k؝�=V!�ٌ�d��^�"�Lmt�85���6F�<��h��;�f�S>����C�Y�Ҟ�q��({��1X�n�����^����S�,�c���6,���E��D�C�a� �zؙp"G==���*A�h^BѬbgڿs�)I@J�c��O�X/Ւ�!��p��t"b,����7�d��g'�����K^ܹ���5n��HSA��hT�B�� �c�J�^���/e�8��!��e�5�`eqI��N���5ȹ}��p��0������0���SF�9���3xTrA)����E5�W)E:�,�V���Ȃ�gp�����2�5Ɨ6ɗK��,�;.�Q�'��Ǩ!uʬ-ƿ&׍\��|Rl�e�u��z�ĻZ���� ��TTE��	�U�j�e��=�W1���XN�N�=������������ȑ,�i�W�9����Z��+V��(X�ǌ��+��`5P����n��쬮��/	T�DJ_٩$��q L��� ���M4����q�(�2��!���x	=�ԓm����BpMf�� �G��
��5}&�兦UJH��{w�.���-�ICS��ގ#')}��ߔ���`I�%t���	��u���ԟ~�<��Oi�k��|�����X���>X
yU�aM�e��+�CO�|�����G4��|�xN��&�zgF���0����]�� z�w��)�/�&�!�KT�v��B��xz����6Jm���'cɭG��;2�HV�����Xp _6Ǿ1����yoo���j�۾�r��	�@v���f�}��n�x8H�n�0�h흯��~G~��R�����g��vM6�9]z^]�x��y%S&�SVadIBpE ����߇VQ_B.K�*ߙ����J���4��=2���}��N��� �M��1���V9f�b��� �#0 ~??�xS�6�I#{-�@�B|~�)���C����C�QvE �}<[+0KP?z�|M;���94�&Ʋ❣3j�����+�2���O.B��A���D��:��l꘣����4���I�@�$��򇥵!!��O ��d�g�=�݈�"���V��:��9��A�Fs=l��0@�����q��5�I$ J��q�xt�����X5���)9��e'E�@	���3ǚհqL������Kr=�+c����P�`��p����3�`�������]�����Mi:}+�ǌ��������V��b0��iKhKN��W���&t�z��
ß�A��ʙZ͂�wt.�/�_mZ���1��0V^�HS�i?Ͻq�$�~�����26���z-�w�;�����VaP:��ZC �H_%�O��cl33�)	G!GO��qk(�g�@���?�H�ޗr�|_Ѡ!�pv�nS�b��'<%�o�����/���|2Gf^��|9��Ux��4m� �̘��3��{�Mh��w����w��֙���ڌ.oئ�i�RT6�>��-��{o#�3�&.˒��8Џc��s�,¬�#5;�>$^� �x'�D������I��g|�f�=]ݓ��h�1��xc�S~ф� .��*���������93�K�9%��z�!����#瓊z�'FA�Qc v�Z�$�I�9%�0�&��g ����qQ�m����D@�a��i��_zB�D@ǩ����I�5qw,�S��"ˮ)F��N�v�m�U�G0�El�Q����b[( �7($�Њ.�FL�4��
�b1��vB ����+;���bo���0؂�5��ǍC���6�)ScT���qhx�j�NH����ho~�>L��
�\t�n.���U�^6�z����	xTE����Y���ŔQ�v��߾<���q@٧0��:��L���#�* rC|��]rJO�R���x�ѡ3�°�&]�4�6R���E>����.a ��K��i0�y���v:�L�`hm�q�/��)��Q�z/����yZ�T�H'��Т���ַ��T�/>K����8'����S-��h#��4���c�j�-�T$���B��[�0޾/[aJIe;�^��8Y�KS^���l���:��^�!i�J�D��a��I2��-�o�M����-�Yx�^�n�*D��A�ܲeX@^dI�?��aT��
���AZɹ��Gsc��.��ٻ@�[�`d��Cw����x�Ίخ�~�ٰI8]����r�����=�i�t�<��l뼰ٿ�^�T���sHD"��k�)����-$����v�#�P�ʽ� yCWԗ�b)��'�B��D�P	��ܝ�� F+!:��
sRb{̡�e�Ǧ���P�-#�̢���%�0@�>Os�>2Nt��NEY�$���V��/
���+����!�&�����~ޯ~!~d���ya*�{0����I��>�
jhs@�m�q����)�Ap�� ?c��Z�4�K�s"�M[N�'"�߹V��/t����B�l�-�U���p��O�u�1 @�b�j���X	?�oK.W��m���TG���5`G�72E'~�/:^������ݿL�=�>��v��Dr*�0�[1�U��A�c�A���E��R��4k����x!&����؂��0�pt��%�LLOx!��?��Z��q��z!���e�ƣ�y՝�/D�-��!�0���~����	��)<�l�+UC3V��Q�?k�M��	$�9g��X�X.h�~�W�/��'��
1��L�{�(�da���^� ��&=��q��OW�X4��V;�Uz�o���WA�iq�"ync8n^t��Y9�
��-��ᯯ�ߋ��#�Q(��^ԩ�1Am��p�|�X�P|E�[Ho��6��i��5��}F�����%;���k�"wC�5"l���9,�e�ǭ��E�З���>b�9�2WS1EI�t��ETiWEI���*������_��1^�+������
��a7�;���
뎔Q�L�A|סI�ݾ]"L˸oOz�	^����'�;�_-�n~3	n�~~G#�������_4��;5$�Z﹍ɤ�T�8�x�ԍs`bH�c�}r&{��=a7Q�7k���J�#	��s=Y��8��?ϭ3n�R �$Ů:��>���or�����?u�����+�̚6xb~�$��0L��E�īcD�5�t���o)��BT\���(�;M׬��%���y��4i�ՠ���qr'��zg*��xI�)��?����X(}T���| YL�+)ȧ�&e�6{ks�m�Rl�3Fe�<��Q����4n��>̯��>5���u�u�����g��Sa��vBSU>���2[��H�	.D.��4�W��Y;i !��#�5�������{�ɑ���a�L����*�b��C+�͚O��?H7�,)p��	����`�p�R=ɞ���N��$�/o��l��ʝ�˹����+�%���{n�Y�##�V`�&qx����:��J+��FKp	�P�cK�~ƣ�{,5OP�~τ��=F����`��Pdܓh�AT�Mn��&A��H��C��Ȯ咏jo�y��RB`},6%b��k�j	fN�_��Ǎ�\F���BLO@��װ6�R�/p�ID��is��T@�/��ǉ
�+�(V9h� �U=��N�x��}���iI�|%��p���Ë��v#��0�M!�zȵqq�4����ը�"�����᳨F`���+�a�<��i�x���������=���A����=sw���C�V�QZ���w����N��1���#Ź�c��Y>���`�$�tE��6:�[m	RzU-i��"��1����k����W�e?��U�$*��.vj37�@���e�.��	3�f����
BR�T]/l]����!P��{j�`K� YS2�t& 
zy�S[Û��6uB��2,��QIf��)����MV��1��ۻ�!�k�X���$�;(&-�v�Of/�ۿ����#���� 4Kӻs���V�|�	6��}2��zv۱�>^¢F�+��Yl��
D�+~D��Ѯ��2&�d�b���v�W����=.F���cc���=:)S�y�o��%��M���u�`ӿo*���%��QΟ�{��.�F���O���s�kU�ѧ�r{��]'>�ÅIIQ>�`#Ʋy���8)6���s��v	j-�l��g!�����_{�@��L+�<Ke�sB��@���l ��U
z�Vrd���G�˝w[k��&9��y����S�ݥ�_Q������畿j�r�F-�Z~A�l��H|c:V�cv� (��ø�ة!���N�T�ة�2r��/)n�j�S����CF��Bt���2YZ�c�F�"l���"��)�_�o����'뭊8��(�>�!M���!�����j!�4Y���┺q$��1��XV��디���>X~x�C��S/�\�I�y.I�U������[s���%Qo�(m��R�}t�mZ?�(����!���'�.H]�g�z�p�#i���\�O[�ǁf���[,��=�.�d-��f���p_�y���A{��X���{���0=x���x��T�(%u��}�}*�;lGXr�N��Ⱥ�l��W�:@���N��i�8�*�PWL�C���$�|�򋳱c[Z�����]�\�yΖ�=����G��@�ߨ�^bD,����_;4yK2�@z��I05�-��#\l�e�?�W����'4")*C^b�j9�.�A-z��)
"��+���K7׏9��㧭l���iyZ�����9ߑ�]�5Q��������ME*?����Cj���Ӕ�۫_�9�n�mVl���"0�/�Z�BO|s�Az��
`��o�2/���@-��Z���M�=����(����6�c���i��D�ܕx��/[�"Ǧ'Ed�TکE\}�W�\�`�k���'o���is��R�4���p>ay�og�"b4��#4�VOJ�k_���+1Л��~;N%g��/��b�]�����Ɩ}���鹘9N���!R��G:>��H޳G_�vE�N���*��V�~��%J� ]�j�z�ʼL����ߕ?�
���d����A��O�w�߱�c��x|���nO�y����7;����5>w8���X��"z�|�'L��w���Oa`P�{]����o�0;2U��~�Y�|�:�;�ɍ��ԣ�kљ�:0��ǳ�qg�J����M��?k���a���G���Ts�q�V���Q�����]�{6�'�u�����,�x���m[�3�^�$��d�)�e�����S��f_iإ�'���"�!Z�Bj����?���$K���O�{H��D�B�y���_@�>ͯ��������ٔ�8���?|�mC�QR�Ӎ竒�'Zp'U�h�l_�h��q�`�U&�eO�����~M�6�kXg/���;�Ѱ��jJ�(�~nG�/��Y�A����sl�g�z.�
�)�Y��c�44��\㮩x3Aڞx"�2�<%|N\������d.�l&�I{
���	�7;:��#*k�b���8���H��$���Mk����QU.�bjn����V�Ͻ��Φ�hp�7��$���`Dλ��A�1�������au�4&��D8<^�&{��N2Ž#:�Qi��ה����)�ؑ�6K��i=��W�ϸ��z�o����GڐU�F���r��iy���s�e�7�I�=z�!�D�t�/�9_�a���+j�#F�3Tv/��¨��C��rJ��hE&{��j�3ݭ�><�$�:Y�<ׂ[[KS�Ϡ�\p>o[�`G���X��I��雨Ŏ�*��=��n��m�{�ד�P�\�:Q*�?��{��f�>%���
��o�va�- �Еg�L���l�U�z�����i�����gpus�Xb��r���_tiar�p
j�]:�*4QD�2�:\mRn
���A�.;	Ws���F��(3��-��	g�Z���3؈�����^V�Q?�E������l,M�sNrv$��J��6dQ37	Un"����|���(n�Xq�7�V�3f�.!|����̨�������1a�]����E���'���_�y�J!c8}�p���>F��k�`d�י �f�?# �w]�ZHu@�&�Sp��0bɲ����Ao���9)�қ�K��|J����XlxVHYEB    fa00    10e0��!u��K�ت���.Ȫ2��b{���ɴ��KDF��|k���R��z0�5տr� l�o�k������GL��-�	�E?n�b�M�?BH'�mE��U<K���_�*#F�n\ZUp���k�L}�s{}�4��	�O�l{ZnUn_��E�\�2��Ѡ�U��F�q�8d
�SCI���.Z� ���ƌG�u�U?XW�뇶�W�V��`��j�%>�_�"��[v7SEg��sC#������};>�c�٬ 9����6i�\�$[���bQ����}.��1Ǔ��t<i}�PLg�j/�|��d��2v�/�*�a�)A�x�&��x� ��kVW~!���V�t{BU���
�m�h�T�YlQ{��)��Ղ�G�@�*d�����Eӯ��N�b�0�qM�R+�V�Iqnkϋ*����jg�\�u��mp
j�=��	�9@�"�"j蘕��>�3_����m�����я���:ۡ�J�����,g�ʤg�-��`�z�Z�u��<��V,��j&:����|�����b)��C�u<���8VF,k��qh��������jM��s?�!��C�����K~��j>��8y�x|T���}TD̉ǐ� �M��g��%�1o�L�G��]��T�[M�i�0����[[e5Ã��Lg�C���F;E�ރHS7��E�}Ȩ}�����$�-�b�|9H��V��ǻ �K���8O;CA����LEl�T�fY-�"M�$;�Ҧc�������,F4���i4MK��*zf����.zު�e>#��&k1���E*����_�ws^��#��`��`����_FYӢ��5�7�Ѳ��3o�qt�p���O:�;�7�����14!)������	�i����fZN
FL@1�s�NY�S���i�n�~A���$���f�8�;�U9��:Uuģ��Y�۬�I�
�Q����ݽX������<��
S�)�צ�"V.R�"�g�4R=�����M�qҨzz�|�{��(NrIK#OJْe��w���d��<�9�����5_�C���YU`A�U�>��h�@�Lx'�P�E��:��������
P�m[�`Vi*.8�^̮`6����$Î�F�S,�@Gm&�\n*5�g�FZ�|�G&���l0Y���ImP:�GxM)tE깖�?~�y�ܖvRANTp����xq�8���m����
�4���{�1O�Q��J��q�/N
)���e0�^��O7��`�| �|��Օ������;F(ς��	hj��"����⣲/(H�0��-�!��:��}��L��z�j��*��Ba���*Fc�x�BU^u�9Pd��E�0���}��`:�j' h��
��w�F����.> M�' ���^8$�i�v"�bFJɎ���vь_����4e���ޡ�~�w4]R�.�r��X��<���9�d`.��-+�[b��x`!�{w�8�5#�݌8��l�2�M�C�����ѷ�9���o��(�(����Jv�=��:!O�ORGF��]pִ����yT��d��ʘ�����=����+9��YfC��Q����Td�,�T3HZ�D�Aik��ٗq�b.��O�|���ρMg�P-X�0�Ȫ��]"+p�l���Zi���r$����c_��+e��8�3)m���t��2"~�:T,K�@�,W�LRLWn�{$BÌjR�]��� ���8o�<Py��'��u�e��P�O���t~V^�]�&|׍`�	f�&�KM\��^�����K+%� ��
j���2#�	�j	朸�mQ?t��ۻO'!�$�B%&r�Ak�p��Ũ�\h��y��U;���6Ua�~oB��K2� ��?�t X�Ɉ��G�do��b�9c۾͵BSh���^�4:y���9! �nH��'�Y*+�����t�t�I������U�!�����'��tL�-Fq��  �'�33ԹT�r�V�]B��ص3C�;.��,(���H�F=(T�!Uȣ{;`��� a�+��
'�������}�űP\i�:��
�+k�5Ր|��b�O|]/��I�.���XV���D����1V���#��4!�V{M�#.�\B��	(�Z4s]4��F�:�}5�Ii����g)a��G��x��v�����x���y8�$�������a���JӊR�G�����ޭ�K�HH��pn/�&F��m������JN2h�A�M*��B ,���O�'>�9����#�&�+���d���Q�g���.B���ë�a ����(k��R9L�\�;�Y�P��E��3�)�wTL��.�]�:���Ji���T�u�͔%(Р�w�&Cg@y�/���Ho�N�x6��k�[�[�B"�\�o�������*9@ ��^ �G77�DP�����o<��~l��ԫ�W����Ӳtb_�Fpy�qz�����[�������{�����>�H1����]}��1I����=&t�QafF�ω&=�"��$p����/ ��.3���kO���]x@[�}%�k�a��?�}g]^�[��8+�yS�8>�B�'O��ٿ�k b=���!�p�[�ia�	��2�o����4�����I��=�"s3J�j��;>
+�+ߐH��fq A0E-�}Ώ��H����#��Z�i��m(Q���%�XpZ}�ɬ�4>;�]�C\��]��;E�-EE՚�*�yL@f�d�k}1͛s����� ���_�����|l9_r�;�H ���d�Íd�S������Ab�&rۊOGb�&�W(�zJ3��ī���6�uzz%��˝ ���D�޹T~��2$��,�.a�%���W��9e��I��w����(".T%��ܐ�6����>����ɓm"�z:-�:���|���;��ԍ!��CA���G���ˍll��D؜�����w�1�M��Ig|�GfWʕ☭�+-�PΕ~I���[��r!	z]ˍ��T�4s�P	ѧ�,k%��řatp�!	1��ڈ�sS�ό�s%�y�tp8Hqm�(l�~^뤩wx+�Y�%W��<H'6*���%5N�~'<T�J�9��ϗ����9��70ʧܒҜ�+ɴฦ,Pv�⨦�nX�_���)�pLE�=>Y��x�k����J"�����)%��d͛��o|[���+����J�qD3�f~�&����F�8�3������V9�����=Rw���1���˴�,�1��G�����X�XFck���O�.�.:�a��7G��/&�Ge?�u7�S�}���+�ڱ��n&& ��"e����XNP�,wJ���Q�,?+�X\�|�\�.46}#��n��F��1B0��cvA��m�[N�p�1�*L�q�p��b�eG�=<�t��U3�F���Q�P��|&������6�92�r܄ѱ�=���=Ap~�1����8�'��P������(��F���h�&³:Q=S:ʲ���D�z�(<2��ĕ)��}ۏ������--�t��-%�1VM;���*6�5r����k�wq0׀�{��i�{���P��R��pJj��������E�~�S#\��
3je��C�rvVЉ��=:�'_!�*Ek��ן�Nʏ�,�k�.8>��ݤr���N��.�f�[5{imFޠP T�(]��9�����-e����@|O@� ,���S|%��U!���^�oD���p%��4-���z����
��j�6�M�Ȍ�!ݮ�.`z:�P0�ʴE�>,��0Jb�����Wi�BU��x��g��Gjӟ�Hs�Æ��s5�[.A�!7���Y#�@�X�|��^��'S�3J6��I\�S����ǡ�Z��&Io�l?���!��B�����dZ�
������x#�X��?�� ��o��������2�v�2�y�:�����0���qmh��ī�~MT\֙J�3ȡ�r����쀰Ta^�ə`%��x�kT��#����_XB��`}G�߫�Q���wi�ٍi_�j�b#cW4�bwϰ0�t�]��E�j~���M ���Y;�+�k�[����P���k4+��1���W��7�I,�Hp��l�aR<�ω�Ss�d�·�&��a	�;����/b��<�[O��]V��Y"ʦ���\Da���v2�_�V��>��_1{h|3�l:�S����f5����3�MoF��� ����dn�xG8̟����iSRS H�����O�XlxVHYEB    fa00    18605�q�k�u�f��5c���Kp�E�.T��V���F�(_�SH@��WR�y�t��#�Q��L���{�f�>�����U �}q�jc��o�������=�Z7W�q��1�@ؔ����3���k0���L�nk��,@��rҔU\�O�8��������W&�~���ͯ׼��*x���l�G�V���@��Y<��8�p���[�du4 ��t3��$�|�B�O�V���AO�����t�kl��d䷇.p_]Z�m 	;U�$
J���W}f�k�ԑ�-���� ���n�8,����6ɤqVE�`�C�SNM~���_�Xx�l+z_W�'ޅ��ǅ�[��r �Ճ��F�Y:?�Cp���)����ΞW�Y��ǩ!.J�2b��6���D]��)@�9��?o۬�jI�d�y�hߠn�o\	x���U���3aG��Q�61�U|��1-����-��գ�����b��˃��~`�I1������<���X�8��t��Z�C��s�RW����<���EW��RB_p�vr��{�[��Y��=$����p��������7�j�N<�s�yt!�(�	,�ª9=���E
N��i��J�.�$��a�x'�=Q��!M�q�U��>: u!�����Ǭ�շ��pٲʐ��8��ֶ���s�g��׀]��Wy5���~�=����'�&���:Ct���6n��7��5�nO�#M9;�M���J�׭�c�)�_6O��qe�늏N_[L�-�ov��X'έi2~P	@�s �iɿǜ�WO�5���&���H����Y�.��Q&KA�=�+��T�9(BoGcb!��B��/N0��T����ѣ�
B��[+��Fo�H�>���1$���M�n�!h�����oK�Ow���6��yض�;��Ec�'��zNa�m�6�M�����AB2��~r���b�ɤ99�@�����v�e�<���h�9�]���^Z���+��[��P}���X�MjԎ�R"��E��<�g�u�j�}uSLS%D���1̦g�M�|��Ws���Pk�JEۡ?�|��l�+vC��I�J��BF9��r��H�a�5��o�
�ߊd9 O�ϸ�7;��NG����2����[�2�t�ߓ��ϑ1��sd�ϯ��0����K�Rpݩ\:,R,�n��Kto�B�nO��, `�tם����g��.�[��j	�ǽ�V`�[�A�*��;K����*��Ɵa�cK���#��L��zi���{�%]��FNJ�ɏASh���0�#�"P�[��S�����e �C?�LhyM������q��'�iW�@�o���S>R���Pt��`T���>�8�^o�+��� ��Ѻ}��r�@Ѳ������*�M�~b�#c�X����.&���|���"�3_S�c�  f9���*�H{�G���v�v �;���f�d� �O-���΀�D��}!n!S��s���2��C��,h�	��K֊��/-�[�ۣ��k6�gy��
�.e���L�����1Vt�9Z�ɟ��Qw,�����P(m�^�2����-���@���g>v���W_z�H?[��A���\M�K��B��3"Kj8�0q��I5a�W�(�����b��-�<��
��5 с@V�8�Hd�Q5r���jlR��a8����[�V=X�I�A�@�Ѣ~��dt���K�Q�=U-6iJ�r��i��e_s�z���&?��J��n�Ac��9��w,�|4]Mp �gu���B���B_��XW��0�=v��ܓ.����`U�DhgE�	pDMWٿ�R���^6ld�J9C��t��1�,���Vfωe�|�n�YOX"ӧN��mFgn%[��(�e�K�����5��%`	��.l@�O�h����GyX�"�����/p��q�0�Mb���F�
}����F�76���KV]G��6�;��� ����D<��a�y��0w���j|Y ���[���"8����E���nL�Z-�b�&�j��Q�cL��4�BY���_�U�պ쓺��t��t�yB�h1&�?�$�1�x)g��&�ϓ��Wb��1��?7Jz �R�\&s��L�Al�3�L���jY�=z����vy�+�����"�$��b^Y��=�ӯ&|sۻfW����Pd��T$wS"��2�	�\~P�A+�g�+��!%͠n��\�X�<+v� ��h�EV�z�+~�Ē�:�+�#1��b��;���.XG�
<�+F�	��)��_І&���o�?Vwr|�H���ڇ����Vs����6��g�ȴ���^\PJ	"ޤ�+���їP�9|�;�C"��3�[�uh���	�� �zD�h%�\D����/�{/����6:i�2�����{��]*�g�i���2�7y��V0!��uQ������YIH��,��n�8O�Ȕ�<YM�9�7?ݙ<P��QW�Nڴ�n ����zo1�Llz����
_	�	���	���$\�'X�8���$�Ƹ����/eE����f��i��x�v�I�o�L^/i�J�1>�>ge˨�EX�J#4���$6<pI��I���@����T�Н��	���z��@����鑹�g�N᧟W�@�y1,�T&3,���B8��u�N�@�l�^8�$	9�n��q�����=�X�@ j��Reo:u����9^��q5��l�;�?Ul��߀�N��Q�������i�P��=�D��WH�ᕓ�T��o�So�����!)��J�10,�
q>X���C�y�.&yŹ��5��<[����I�k�i�������V6��o�j$���k;,1�e�t�(<��[�z9�b:�3�[W�U�t<l���淹��*2C�_��$�[�4Għ��Et�~n�ծ� �$��Y�K
S�"��WiD��F��k����퐢���E(���ꨶ�"�p�8��|Jɹ�j��\'	`ϐlkZu���KBv�P�/����Ux��E�8G���u�|��(��~��y��g�[�g�FRic���(�J
>63	B@�IE8�ı�O�*�PS��>*}�l2Ӣ�.���A$�	�am@$oJ��F�K���tP
pg@�g��TSļ��M�C1>�,DѕFl�x7��FC��^�#�.0*x{��'z���f�f{>�Q8A?���E�ӂd�V �n��V���j����`�/K6]�5B;ꑑ �����b�� �t��"�X�S�����}���� ۨ���&�~�ڰ�1|�鰡l��/5}o�''E�X�,�{Pl��GE�� ~4�FAyb���M���Z��$ >:2�v�M��4g)r6o��C�2����nZ�A>��{7#�2�Y8��:Ϩ��K�e�O�WM9��x�gk|o"�Q����N��,�<QG8qZԷ�{�
������p�[��m.�	�ڬ^������6�����B������x��w�]k��9;�,'Z�*�W��`D֛��d?����d!��莌�-1'��-��y�P�ǶA: W��6�y.,[߆ д��Uz�Wء���>d63��8��юJ��$O�̇�y�/�q�#+����u�#���/��).�i}	��|��D�*Z��)yB� �]�T�^���|1��A��i��6�Ώ�XÃ�x�e*K�>�Ҩ1��x޵/J�l�5�5I	W �+�
QK��T����gW���[��>��fB�jc�������`�|#���_��L2*��_�C�M�2�|�Z^��X��#�LO��J��t ?�S���yU)�P�aV`�Ϝ�s�a"�?{g�V�&��P��*w؞�E��L������=�����%g�6&B>��K���_z|�u���8	�=^��)93k�ۺS"+�3��Pٰ_�T 2u�C7�1���-��"��S�#�63n/�x>R{-��3ǢZǏ�����dj�� �0��!��s��]I��x�ߛ`�Sx�N�����3���kE��1����ՅF.�&�i�i�R��G����7<�D��Z�x6�1��\ k���		�����W��(zQ2��l����%O�x�{�]�� =eM�u
�-++�eSn;������ݱU����v�w,n�;���C7�s�*t1��H��gz���<�j͎1�q~�E�%	����l���h�\0��z0b҈�&�������s��>�m>�૳�o߬��v����2��W)u��x��t���Ѩ3����f?m?�U�����D���2�|��[pp�C���h���:.�p���uG�,���)VQE�T�+�*�D�v��޴w�?�� N�1�=�+����8��f�����/��9N��v��Ԓd&V��kP�';]j���jLɹ
��'�C�ƶS@��UPq1Z ��s`k�P��ZiU��j�����6�@4�U���ߓ�gg�-�x��0o�t "@i�#Q������,�č��y�h@�1e*�|��X`|�>�p�jcWQ`)��9�}����w��\lcu��sT�OIBr�q�8J���R�f�vR^��9��Bo�;E��ě���8��)�9�Aa�ƍ��C����V�%:54��Ԫ�K� �b����'�+�W=�ܷ�d �A��	R���2�: �7��*fʒנ�� l8v�5's�f�?�b��˫���*�!��d�ǽm���`�a���wW!�jsk������:�Y<ɷ����a�F��1I>/S��]�z��QB�aQ^�ALU��䭭�CA��Y�9$xد���u �tu��sO�BX���j���W��pn���݄��0��L���P"�ë'u��ԍb���<�99���� I-���an�QkO�L:|��d��m��G��p]Q<�Xw�^ۗZ�z�Eh?з'3��t4��� �U�6W�Q������W�ͅ�\ש�Q��;�����OquLCy�����|g�;��0�
s�>Z���(^<mp���Vx�o��[����Y�dGK�[��/�n�i��7��d��o�;�0�a���2��N�xIkr�j�8���J"���s�&wMMD��p�������@���2F�Z��<��&r���f���V�PG�.G����IB�S��Lj�����n*��]F�B�/,���:gXY�Í.XʩY�b����ެ�0�M? �k���4t2reqeʈ��c��. jC7�p��.��m�R���L ��������A~���uY
�f�Ş~���t)l����$�/+�#�Pvy�~;���do�;���M����&a_(�9jSM��s��VKg^1��2�y�IlTY��ƓM���S^w��[��JuI%_B��� vW�x3/��X �;R"�3�(���{�=dmW(���N\�f�i�����s��6@� �,��Q=�R��9q�7�æ��
�\�:����t$�2 ��T�nh�����6�4&7��[�f3h82Q$;<ܞ��Y��u��Ӕ�[�_�U����S/���H�G��]�o�}6��f�͋�n|>]ݨ��1�n�֐�͹'0q��� _�෾)��C:&�����ZH����K��2�~�E�^���Y��9u�,fa��W��xWЌ�Ґ��GN���C���ץ�O�8u+�Ez~l��d[O�ū��.`('�NW⼤��g��]B�ؤfF��Эc�h����/�y	 P���������ue���ӥ'����N��
1fg-Q�=*i���i��P$���I(a��[E����.�0�ց:��jy���*�̒�H	x������6�#��I�R÷Q:�u}�nZ�O���9�0(rI�I[nLj ��G��ݼ����)�g�ʐv�����^�ak"D*��4��1#۰�mͿ���B�/mx�%�n� ���'��5��i����/T%��+��7?��zOO��x=���|�"�9O�%�E����"�3����c����*�4�55�{�o3	�}��.�O��L��P�I]��xw\���P����|^5$MS�J��qU�jq�{�ٹ����a6ng|I������u��D:Y8:���f�dBY,w��S�,ё��TXlxVHYEB    fa00    1720��k;�X� ��'���i��|���? ��J�SY6��ϼ�A�[�dI��w�fk�)�8Q���f�p�ߦa"*��,�W�u�I7�D`�~�X���q��Uu�����3�t�^�z���z��ܡ?�^�`�;i�0 �,m�
�*iɣP�CHH��V-���K[Ҳ����������Ik >�3�����T8�n��#$bw@��*l2<�RxA���A��֚��ơp����`����s~��V�r�Zo��xd��6'o�'
�GS�4=���h�xM(R�rD]N߬,ӻ��sL�ڰ@���y�/Y:y��8�>��M���:`�y="�Oτ��EO�8Q묶_�H"r���*_�RMd��b�iD{���|��|��|��g�mP�๢���]��8��jq�(��t�eſ!���[,�p(�8���\(k�-��Ʋ���w7I�ރ'����yy�|�-���d	/��5ʁ������Y�$(���>ߝW;,�����t���o����O��C
�#]QG/�[�9z +�_|��fTy�i2�N��⺵M�]԰JI�k�x�-{~K,jb�կ{�§����ҥe(,���'ML�c��1��C��Ν�ՙ�hla�#JI,�d.�wʱg\.�\���ku�n��+��7�˜�ӑǦ��5<��׺u��� �zR���h6��D��:c��S5� ���1�?UݶJ.i"�_I�+�w{'�R�QFB��a;!�O6���0�ԣ��������B\�^�򛋉�d�����/C�\�VE�x4�' ��x��D�^�g��h���\�r�+�7i�wbm�Bγ�����W��c ��u�;��04��S.���v ���3]�%l�*?��;��)�뮴�������r�_��}Y����D7�Q~X���Z��x���R��7���z�����C���nR������{@��b� b%vG�-j�3�)��C��� ��X��2E98�%bA���Vo�ſ�c\�8A�	i��&�����h];�6���.6H*� �0�!�.WE 
��-ș�Ȼ��Z�y��I⬉����sA>�#PV��������^�ȩ����2�׼dy�����y�@�2x/����)��r��mm @�VYI�o�
��>��s
��E!���W�'��<���/����i���h���n�X���;yFܾ�C��႘%N��MϠ��2�����>?��|��`��z����d_�������V�|aκ�5��ȭ}|�mjq�x����0�a[�՛�!��~e|�ָ虔�g�h�	b��H'0���{[�5\e�]aL֡3�>TO��n�/m��Ky�g� �a���}�.�x�����ߟg�'�����J)�}K����!aXY�sF�GA�;58b^G�M������
��*8ҹ�m���w~/;�u�vWw�^���!$_�|0���*���4�B�� ;��y���:~:LsQQ!cý�����mW����;]������N�Kv!�n�{`�ao���>ˑ��1	����VQ^A{Ќ�!L�<:����-M�P�i$z�u��V��ۚ�e$��D&��S4b��XÌt����z:t���V߂?�ɇ'�������.kmKOENf����b�[+������}��!k5�S�,}�I$��i'o����:8�� ��z�Kƣ&\k^�j1����MuKYu&�֥_�=\��s��D�7P��o9L�٠��&�L��ݩ>{�3��2�;��{���!K�P���JXL����P�1d�,�q�Q���_;<#���6����~��������?y��R���Q m��$I������QJ}�=T ҋ:�+!��/l
h"���?��q6�u|�O�ldS�.%��lc����>=N�y��Q���v�U,�V)z�k9IQs�"v��n�����e����W�3��?� �f<ݯ�G�}_ϰ��&�]/�w�~q�޻�gH���o��>8.Ұ��,�V?�N) �-��"#$]V�u%t�6�Ϣ���^[c�3�S��P�Ӏ0w#��V^�ӊ�z�=�S&/vC8j��'5/��

���J��8�3o����#BT�K�լ�.���m@i(�A*������a��s��uo,����L��?~V�ϴL����}y$ױh8�qd��B,�����2����O�94L�}��q�h dA,hSH[8�f��>:��/�%*�5Դ욟jQɓ'���3���$iO�'H�y^�-t)N��6�]��=A���=b�\h��+�V[nC�c�W���lY����Kc=��)Vm�
a����إH>�.�r{ZP��0m�|���5�-�<Ż�l4�Uo��g�0,L��(U���������ʭ�3y���~�.ED�8��2�['�Z�-���V1�	�F0f붋��J4�� 7e�{��7O!���qۖ����+�4k�'�khfEX�%A��9�]�����s<޲�ׯ�C��3W��B��imx��՘��Y̐,��%��4�r�QhW��H՚O�D�����4o����`,6!��i��Ǵ�~��ݥ�O��V�*[d�W�o|~��tu�@ ���x]�I�ad�0��@�?s��ɗ����u��<�
y��0Y��@5woẂ˂��Z9-M"{��)]��-�n(���z�5Z\tk�쏌{��k�f�``��G�]-%��g��@��Yt����Ef/D���,��2��{�������:�:'N��6�8�_V?4��K�փp�9��_�A�
��krX����N���|b�le*��넟�ό2�&�����ܓ썬��Ϸ���8��n��
+�!wVT�|�c���H+A�*y����Y�y�7$�vC6-\�t׼��/6�O��� �"�(�m��3�vL�3��ۅx5�X��*��1�ь�?K�'�+���H��q�����%��#�r�"������I{^�����Q1���;۟��n╶��!���P���*�;��b��w��`�'���A�j��ﯭq�C�^�:qD�q�R'jh�CGJ�^}�f��*Jͨ=0������!q���6� �1�LL��^��6�ˉH��QB/��VW����u�������>�&���OM\��)lk2�Z2���ƃ/�����!�l߫�&Z��Fq[�b\>c�eҏ�+��j-m,�����7�з�,�#�MF*s��9�#Ș��r�n���w����Zo1�3�'��\s��;6�3�`���B~Y�uV�r
��0�?������\M��a?�����5u����[T�m	��%V	f@����0�7p���ԫ�B�0�)�I��\�ȧ��Rc���i���>,��w<��h��HT���t����DcATW��]��3�X9.F�ފxK�+=���Y�(L�ϒI< ��� �f5����"������w^��Hz4K~a�rQ	�1�X�Ub{j�L|��~Ϗl�bL�7��Dd�TsJ�^܏E�U�����z2��w�
OK�o���ԗ��BPB���zZI"�l8f�E��Z��	�|c�W�"Dt=����k��<��(f���C�&P��G棌�������u"�Ν����63��pR�<����m���q�����@y$����:��L��Ou��>�~��2��Mʮ�90��(=�Y=>q��� �m���V�l8�Vd�����m�􆘰�;vb�l�@JY��p��ڛ.)������Mմ�Iz��y \�-05N�N��q�9Xu�� ��ދ�������-�BnaQ��лҍ����U����ϭ�AX���U�q�)%UH������GKz��S���\�����l�C�@~�!�gw�o�9��l��3kp������G����n��aI�_$r��s40]�^�źBp������['څ�������:��(����ʒ
A9�U�&���Tw�D�)�<�-�q�g�H�[B�X�	�A�ܷ<;k�ٳB&#K�I2w���v�~=t�\�z44�k[��J/��၄W7ȿ�ˠܣ`8�fٌ;��5d��Jjc�t�\a\l7�� pul]8�G(�B�>w� Oj7�ʩ��]��	kzgQ%,���r��ݐ;@�{K%���nk.�:%�����<�&JZp<κr/���kx�b�n!���vŖ�(K��7��\�ȕ���=�SW�2�&�z�;1P�o1����~�sm4O��BG���R��(��K̉�^+������6s�=sa��j	j����#Уs�ݩ�6�BY^�%{|r�6�oW�*n���d����P"��6A֣����(�&�!;=Z+�a^�'�M�	ފuW�{ ���������I�R�o�.��25W�Ԓ���xYB��������ac:����I6�[���H�b�t�35y�(�Y�#���ǯ(埥(�Y�v�s����4n��j⪱u)6u����B���X��Ù���z�#2��U
\�-ϩ;t�S" ��"�M��K�q�t O���S{TG��q+(�	4;1CR^�/̆P*��Q/`��0�Z��A������БqY5Q,���͞�9��Y��2�,ue��}�XGc �o�O�Y��Bd̵
Iן�ǋP����Z>����'�;�69���*"�ͣ�:m��T 3�}z8Ơ���B�R@�I����O�;�71�<�!�����������1'�T:��Q�mV-��/��94�t���upī!1F.�WH�ֻ<ulJ�
�v�y�茹� ���ʀ*s	�I�'�aT�ZR�D�it'�J`�_`sTu�����$-Q�EP>���D���+d�x�zpK�*�
ぃ��4��Rw�x�Ƀ(+����$��7�tp�
q�
���W`a�s��c��I^J�E�p�=�6��S�j(���p�G�������2u!�F��.�O��J$�j&���H�t�6k�йU���.�3�	&pJ��1�MU��x̥.�	^��c��c1�a�ݺb��o�2*�v�����
��uQZ�e��a��t(�	WFt�NS�DjТ���>��Q���5�.��
��6\h8���a^2�r�M���d�g�%��'<S��w
k�<�CL6j�K&_G��,\e�
���F5|5n��~^�&���E�J�kTv�/9h�-�u��'�P��|�s��=s����&˦�I�[�Se��@f� �=��2B���ZW����&ʉw�E��s�$��̺jǀ	z�n�#����j9�|�, ��7����0i���\m����oЕ���(�4y�r���>�c���(j�8�Z0�����q�=C�|��XR@W�C�Հ';<�v�c(��� ��6�<�k�1���B{<�Kl�F�c��:����m')��ay_��Aa�;���G+𢬠�c���	Пg_w�b0ĒQ��K�x�����E	���TR���(6����@a�^Ms�.���L�f3Z�M�c�(_�B/�oE�i㵵*t�.��kH��1�����i����	�4$�<a0�ok@�����z�.3�:ם0���b9%z�4��Ƌ����7�M�9X"â�6I�܎�S�li�4�)�^��Ip�c�-9~���	�F�G��J��$����\�U̫�j�}2����.Ii�F�s2�Z�r4�D;Ji�T]�@�r�<Y^�����?�ovHA���8��(wG��'���f�χz�d5yٺ?�]Trق�rN��ylasў�p�9���%s~�5yuR���n{��PCD��mr��ѵ�X�_Q�/?˰��¯$�+wj�mĒ�p����h���'�I�N�At2CH��1��W�7�!��XlxVHYEB    fa00    1500}�ߌ�M�j���K��pC�ϣ6<�oZ��7��e�_
�	�W�4k"����t.Ø�+QY(8b�q6���J;��7��o;�DL�#��уNC?�kC�ڥ�#<:Xĕ�A�Z*���
+,X�C��[����*a��Fմ\�qÈR���
+�����"3��ɢ��~��~�v.Y9���~%<�Y�������/����	P�:J~��;��5���g\�\WN��"|�F�B���/�)��Z��A�|wC�Գn�t�C~{<��R!���ExS�����H��i`� X���԰28�T=�U,FL3O����A9Ou_�4����DJ���!U�3i���Ǚ��U_��^a	fF��U���;��̈�0�_��v�	�#��zo �2N�M|�py�^���U���lƷ�"3�4�����.v��։6�*�A���]v4`#q�;��Y��i�����m���&&t��� L"�98TK_��*��;��ɐ�}`�G\�XC9��4���y͞�s8>�Y�ʰ_�k�2��]��ӱ�V��BxY�|2��Z�ݕ��Ӫ�zDl�Y���%ږ�5��%`Lȅ{_�b5��h���{ws���/Y$⮃�M�ܭo�,#{�6q�]ɲMm:�:�J�[���b-F���Cp
��H��b��w�m�����y�;�&�ƌ#�X`�ɖ�Fv�.����! ^\وH[��p82���j����U;��5¾Ns�h���T�W8mF��۵`R�$�� A[�V�7���(�1 V��F�۳��h�'}m���Vi��+��� J��k���e�)���3ie�j����>���Y	��{U���rh�/��)U�j���Ga&	��q]���"��Sp�G��� M��0W��e���ۍS#�1J��S���-y���mܕ!�o�Lw@U�2:ߝv�Φ�7�l����{�kci\�-b^���j�s/Ax˨�%V��Ϡ� e\����a���<��k�1B��)I9�(�.��8|�+	\x��Ԕ�rF��߳��!��D)U�5�	m���e�u�B�G�����\M�`Zۡ�1�`f�REi�߉hAf�Ц�n6 3敌���g�u�E� �Q�j��3����FPf�A���=G�x�O+c��![5a�%�Q��]�uu��&�>�P�b�I3�Opc�-RO��Q���X�j��<P�S��~b�$Ӈ��/�!..�Q�Sc4�#T�qB�HB��;��%�N%�f�;�a�q �\q#s���9ȑXgs/B�5߃XTg$����b����Y "y�Һ�-���j=����HDZ&��	��Uhwͫ�,������N���2���&9/��0��*�G�Q��w���~ԗ̓7a��w	�ƞ����֟2i�iGA�%��ݾLp ��Fg��ƿ��ă`�=
�4�����r.v���А�(H���{9 �SXY����#�z�~�}�W�9���.)5K���L�J�#��LP�@�D��-}���~K=.ˣ��J<�acr�dI���>`�º��ط����� �m_n�P�9S���5^�\�j?�ptvs�l\t�1E>�c]	\��EI��/፵FfxD����7�#�_V�,�&���QLn0�R�ƽ�`�pA�YY+8��u�{#���H�z�jw�<�L�;@9xk7@�FH� �p\�j�M�A@L�������W�AU��Fޒ~|ҩ�<������U����J<=�%"�R�&�x�I�F0F/����1&�,�f�8�Ej<)��K�6�AÔJ�1Y��c�r>��-M��)v��I|�+o�ו��?�R>��q*M�P0��'X���1�������@�����u����M��ƛ�����1��~�_��֘f�0��������4�g�<�F�J���gz�X�Kj���3��L*J_��"(�j������_-�=܏=�?�{I����}�W�o	�ܿ=��&t,o|���O��MV^����Ix��B�H̏��W���*�T��ZN��eU��Z�`�˨6��'}�����!�����se<�Ӊ~� y���Z5;r,����w�A�澗�6���]��0"�w�����9�V�����0�U�)aw6��c� 3R����é�����/ȅ/~��|>���k�c�Q��&&m��:]%ɓ>*�,����[�+ZOo��"���[Ң�����ˬ�z�h4;�b�U �/�/z�\*���P"���qo84�e�6r���{X�8zǁu�0z��q�,�LNDߖ��.���*.��v��!��q*�8��IkD��~��;�~�����%�N��RQ��Ė�r��n�3���8���ʧ�V��;Q`�5�����3/AOO�����|3�ꝀH�gv�Ẅd���<�{:�w��Ð���O䔃�����gVi� 5�S�2ԄHunl	E�Z���~�ZLG��iP��Q�B�o�Jt,�Km��PQ��l�_�
nZ!k
�/#�T�h�
��&`+@�����yoY�S�p,�%Q�����Q�3`��j;�T��lX�PJ�6���x:��^7;�[ߪa�9��Z�L�s��O�R�+!��c�dD_�$;k�⁲x�D���E�R��N��	�C�#f*�^����/~>���p�Q�U�-�2H�A�N�`V=0^��[cd��Ɋ4��+�m�]�Y�ʌ{�"������2r�P�����nu�,�«ONuI�Ppa6����<��2�T�w��L��YX�	�u��jǆ��Ÿl��}�M5�d����f���q�&Z��h�߈�i+i��#s���y��v�k��[_���T�y��щ���h�[a����50kΗva%1�rA#�E)��;衞�����mf_���H���B�-�i	hD������<���
,��oO�MpZ!%�H�'c]�ϑ�~k]ׯ� ���{�Cbܾ���b2���R3C$4>�b@n�'wA$�\�M�ȿ��W��kH�;����a�~�R�ڻ�7R��(�$�m�ȟy�)Qk��[D�^GO~�����	m�ŗFu|��V
��)ҫ�kAy�BՏ���Z`��l0�[c��Hw������<OJ�D=K�/�[&�A@S����rePNO��:�I�tA[��6$�d6	R��p�1�j�����',�x�:A�35����U�/o�J�}VX���2�ajF��X�q�[jc�8�O*-��y h��G�T��I�?/ff9�����}���y����;Z9Z�0c���R��Yc9��?=&��BK��Sӱ���,�H�]�~�$��[P$^XU�GM�%���ɠi.������ތm�UD�d={��uM�s�ݴ�+�-�(��	͔�.�{e��3�ǹ�?i���K��/��׵[���}�v��� ���`e[i扫�2���r��QbM�fԺ݄�;c�}��� K~��_-�%�>�e��=��-fiy��(H�������~��8:_�
%QD"�$���O�^r^�yF[ǰ�t�e��K^|��j���4Y�7����P��Eg�̫'�.2�?�+�(�C�A3l�#���%��z�QG�W��^�S����	�/���p�+�ƶ���h�\fJ/gȀE��B���K�zs���g�TU���-�b����P��b�K,PUF"Z
7m�JB�9z����T���v�R[�,%�Q���*&�/��ç*��O����Ѹ(w���? 1Pr��8C=���XwA��,Ɇ#����N���+m$�-��0)EM����qa�Gw��O�w'���p!~��F���G�9��e���Ʉ����N��XEuj���'t/�|ī1I�vI`�_O����	x�r�f�����$��I�������d}'�=�# S�]B�$�o���b>v��t�f����qeԘMY
� m��5e��hz?߷ן��Պz�0!����!x�y�v���,]*��!�N�l1Ws<�D~Y*�\���b��2v�y��nHK:IK@�^a�Ѱ��B1��V�-���Y��y�+�R<dI�$%�4;=�^�X��#V�L��sP�2Ơ|�!�vu��`�5�Kf0C�m$��|��BR-1�i��{5z��JJ �!Zv��ʲ(��K��f1�u����oKx�ۄv+֗���0����O�6�ؤ�l=�0��X8���Νz~�i��D��	�K��,�
9t�Tf�3���X��Rq8-{H��t���Q�w\��2�닿�g�0��=���)�V* *-ε�F��7��u ~��dK�/����6��<Ȥ��	�1�]�HBB�a/z�U0�J�)�K7WO��޶1C&l���Qq�jX3�������Dd
'O�?�H�� d�+I��;��H��+r��xb�3�R�L%)�'�]��]o,AT�N�[����g(�_^_<G�uP�C�TG��/o�P�|Ǫ�,(������ي FƁ��媉b���ә^�B�:K�e���s�힊�m��ZL� �=���0\�3Lc�H筠��;���$5��p"��|Qp��U��i?M��P�O˻��S����#-�G�'�r�pG�xw�j�j�HC�4�^Hvi���o>�u��j�fd`��쥉c�We�IH�P��r���us��æ�$}k'�5���.bM��r��U4�|�8�gmP���}?a�}Ľ���
S0d�	#0dtauij�S���T�f��KK1��}�nsNf��h���?����n车hv�o7#��r�˘n�[ȵ~���hXC�t٦3�z�o��#� ��E" Q)[��G@E�A˵;�ϱ���w�)!�wz�~)��q��n�ΰ�x���M��S@I��H}�ș�W��!�ۢv{�M��-�Շ��:H겣�,ȑ>��o��`§�K����MƟ�Q&�k��Q�?c�|I6_P4|%k��.��D�Oh��4G�"�iC�R��.y$���y��4��>{,�Vo�5(�=E '�X�A��%�j��b���!�@�Za=�P[�_�lEЯ��{�S���1����YzXH�~�$u�$���֋Yb[u�*X]�0��&je�*���X�����e�����\�9�c�6���cqGTl���l���
�6I}+�՗����CZ�kLC��*����0��=�b���*=�^©|��c����r��������9�P2�Z��}z5>�|Q/���xH��o^�[�ߝ�&��>� [;s�N8H����E��| t�Wj=������>�C��O�Ŵ9�06t��XlxVHYEB    fa00    16c0���InD�%������&j{c���~W�:O-�3@��Þ�yD�X�o�B!m	R���AcS�U�UI�Q����6�{lХP��K͖�٧�+K���]����%j5�A^���G���K�&�L_lSV�6�p�dB1{M{=�7(a��H��}�OLw�Ÿ`P��}H8�.�\�<G,B���Y���䲗-V1eM�#Ѫ75aF����E��;��ݩ� �������
��;�Ynb��DQz6Jw��3�a�-ɇ�����y�ţ8AE�4
�}���	�T��b�}� �X(e��*���4!)���<	�_"�	y��%`��R��ǌ) &j��~����.��F\>��62�����{��*�mH9�]fv��F'�g㄄"F\i1��z��&~wk�;�<�),��v��5�p-�Sg�6�P�ɬ���;��V�(�m}#!�k�ȸ\��8�,�
�Bw?�*�=o�%��a���Aw��ڢ� ��������qQ�P�_�M|dhHD}�#�t��R��p���d7W���ǲq���,c���I`ֶ���7�~D��Ŭ_���%���ώ̨C�"$��f$Q�7���}������x�MA�Uy̦T�HB����b�3�w'����I~��ڍNﳣR��9:�R�Ț��tp|�c��"`��Oq�kVʹ�'F	���N�	h�Z	h�B�F�z���^D�g7��Bɐ6y�z�IZH"o��[Y0}4H��t��A?K<O�L� ��~r9`vOJ9�s�r�n�J�BX[X��\��F�<H`�:x{�y���.Ib��D�pW�4䗭U��D؃-�h�Xꊼ��k\g��0�#���.V�r�s����4�;���N��}����|�#o�#��I3Y>��yx
��~":_.��pRx9[Q2/�8�M�]U��ѶSN�S4�nP�2���XL��E���b.�TݷU���6����>�}x����\k��o��=�
�b�z��"�:��?!qm�\�s�L�H�9��Q���^���)kQ.a�o�譄ߐ����Ped["p~[`l�b878y9��)=ퟬ�2C~�������R���7��(l��<o���ʣ�%t��%��#��K�fO��e%��ܷ��?I3^��s��p��]����~�"�O�|�"*v�'�9d.j����Z��AB��߷6{]o�*^��,\�c��![2)
аsU��)�_�ik�dH��b3"�_��,���&lb1�7�-��(h譮����ߜ���u��X}��3f_4�]Qq�j5�>iJ��J1�QuL������|��a╖��Dׅ�.����A�/{>�|b/�W NOw�Fl1�q]hO������($"��c�&��@��*���kXx�4Z�w�.��^�TF�%�Ad��xX��kI ,�/oBw�¦X��O�]��WG��Uox�gtkh����c���xn}>���!X
���\gS$S8L��yADZ<bJ���E7�j�#҈r��|(0����Gҥ��(�Bi�8-oc��e	�JH\�=kˑI�:���i�(���q��1��I��ݦ����D������$SkFv;���&=:�W��(�� Gݹ�-���m�!j��MА����A!N���3г�B�q���p��o�P�t�Iu.Wـu�V���K�#��C�*Zk6!�ݖ�-�����3&$c�d�qA��X�F2�,I�좂��à�T3������TќB���psm�o��v��{���3�'"� �a�Ah��^�Bv�F�+G�w��Z�7��4��o2��_�k�y��1��U-��"�ƴ�v��D�UI�E��?�	�$a�k=��m���tJ����G�����y�;���f�� �J�[?�SNT_m�cYn����๩3X�h�T����؏J��.iN">J�%�$��Ӵ�����ѥ�B2���!��� =��<ߙ��Y�	6��L�	w�+
nz0"%��P���i�mmt��׍Ib�}��u�/V��.ǥ�i���d�VwV�2t�B_��P����9@�:���cp<���cZ�
,fO�n�����{��6菕>�&����tMPĬ=9NE�]
ᓣI]�"���u��fd�!W��},`��jO�<�u�:�Z���*|��&(�ܜ��*�P��'����Db�Pi�~!��|^�cM����[�|���!}g� <���C����{�2RRdÄE�80&�ٴ>�9�z�SK�o���[G������n�m�0$�`Qp�I�����Ҧ'�'�^d�^(��t6ӗ�����f��������]3x�;sS|$2`�D_��^���BU�:�NO��n%Y�P3O�L$��9�K�8�6^�/tt,�n������>$�۲e���U�l�ep�E�$�G�"yA�he�A�Q�K=���
^��f��n��i���[�h'��$�O���竛o4����It��LI�oMuGMg<ͳ'��(RD�<ǝh+:W���MKe���(쬃)����Q���x$P�O;�]��s/��(FpS�`�W�M�O��9�ԯ�����ܧ�z����,�-�z��}�"�x��S�#Bƣ�֍K��O�I�ܝT�zr��C����2�_��>�6[�;P��]��n��j�)��FM�j&o<O6������<M�>�e��TQ��d5�~�N�����+c|>@�謰�����R^ �h>������*�V�H���ۤ�.nȴƼ���3�ϙaB����Og�ݙ���𶧾�43���n粸ad\@� ���0���.EB(x��),�S�[y+3q���/+�����elI�m2�����ط�b_o�F���>�XwZ�ή�t�&nrșK%���92k|�i�:�K���9%�Ց���P+�F6��+�ȳ_�\#z��Z|@&�Xէ�X��%P�JU��;�}�7nPx��'�ݚ߈��������8�����s�?�,�Mc�<5}�%�R���#��h�#L�>7�4�����;^^M/��\~|0��hn�)�i�U��N͆촛�=�kՔ$���]x�O���/1F ��
@t���Y��Æq������.�|Fs��|��$��h����S,zn�����^��?�����`�~cf#eE�{��՛�����5z2z��I	T+
�k���!'�*�P��Ԍ������"�C���؞�[��pe��[w�9������r%�}�\@�D W{��5&t�'���$w�&�oVJ��;9�Ŕ��Tp2�^�?��F����.�6�{�W�O.��EB�C�Y��G˱������ �i��1�Q�w�a~�!NF�@�ۏ�s6�T(m�&�!O��a���V�gy�Su��7u�9�0�3��$A�]4� 7��7���./���؜�=�<l�F�ՏtOu��XK� ��c����
)�8�;IMEw����|���ݸJ;��������R�\8Q��8�Нҍ|3�|��:Z�K��ח�{�-�P��lS�XGl�E����uZ`��%�2;x28UE���pB�{�:̤z�[�-��'B��;�*y\���k��M��tBe@���y�N<KK#y�Uw�!;h�A�����Gm�w}1O�E���#n��V�~u�m|Np�CU��;��Y@����쎔�+��X�ʥ�C��5Pw v�����o�L��r�kA�&pq�����o���-�Z�S��;	�V2���QA~�P�_��)��A{��1��ʎ�S�Yu֊��|����
+�O���������
R�x*�>i�W"N�d:��Y�H��o��3�|� �M!g;dzs�܀W���1�M^˨�@5�l�{�@5��-D�M�vus!�m�-E�4c������0]�&��$|�����&�4XH�p`&#Ѣ@}�3�����f��̵ؑ�E�D�nP<q5��ֈkИ4��l���t��I�{TU�r�� ��{A/��z��VZ��S�汻{-��b�����8Q?�eCP]�����79�	h�Φ(���E��5r�g-E̗���)���b"���1��j��Z��BꞈNta�C,�$�4���p�Iܽ�xo+��K'���
�TL�%�j�|EW
���6�'�:�������&�5�q�V�G�gk�H�5l��/0�a��TG���8u�2��0��O~?�+ ��j���[�kd |p�-�:U2����1���q��ي��E��:`�0A��rq��C*�_�q�xaT�wM
{?�U����>�l��	T_��;�t�B�Y-��ͩ|����x��$�
�3Ԍh����qCw�$�>�x��>���~�0	����T�,�'�<9�qՀuC���k%�c�p�{$o�$��qΓ��I|��Y��� �6ĵ,A��|��zU���� �Z�_I��pt��5(!�@�i�S�1�I���w'`��G��Ux@1���&�?��E�'�K�r=ab;��<��]��dum��Z�pb�F�������S8��r�2w���dY��8 �R%�������.�^���7�,����K��O#j�a�+�w;B4� �|�UP��(����ܯ�V�V�wq���sd�&��Zx+{�����p�L�{}�2�j�-��oy��ʯE~���!��k�"l��6�2�S!2�,�����@��ސWΩگ�;H#ղ����f�n����鎪�e�Z�����Qxn`X��C,�rB��gx3:�/�U�M��.s��U��8�|,��]؄���L"X�EMs-+����{�p��0�^eԅ�ꫦ������B��`H&J�P_ͩ4�-䏓)��M�8�L�?�:�y�R ���KQ�	m��F?���=�Me���X%/�Uʹ/f��
z^"�~Zn��IƂ[�n��������"[�@�g��o��b �H���W����Vde��ySi��<�D���݄�C��<��' �]��3=
�z�m_P:�/���e�z���5�(�u���WB����sCӋWD�������<`���U���B!H.9d)>�B+�����o�)T�@(̨��3���M�f(�N��"���wH44�� H4�ۄh�{8AB�sY��o(�P'#�@ �pV�>�B�@Xg��㮣�u�e�a�'�QS�s;�F,���&�2 k�rׄPlf[X�X7���F���B6(�����A�eE��ј"ȭ�X�'�2L�/�Y��x�q 's�̃K,�M=�N�>��C��!�E��כ3�Ex ��øWr�Y�����O�5.�-�>��>�T�1�b.Z���Z�+ �)�R��%~7`��]4Y&��]��d�Z�����9�0�c��VZ+�,�V]e��xtd��I��و��(�w{����ECn��Ev)\NS��<�����G����
g����-V�b�7���;BpˮBo[�۵��Y����A��?���|����T}�?��tҳqAf�!�Kv�L��*='T��1��~�P�g]��uIy�Z�"�<s�ˑ�嶒�t,�cn��t��}�4�Dur
(Tqe{�����I�I�F���5�X���f~�|�n���\�
K�/%�����Y3����f���G��%s��\'\)w;ݖ娃\o���=�V �"X��q��?��F��q�ڌ
hV^�q;�� �j&rhj�7��LyŔ���M�2�N�K+3/�ʽ�Y9xG��rbXlxVHYEB    fa00    1740!Z���r%K�p�`�'��YHfL�-B��Z���L~��R#+v�?�|�PC�<�4�W\?(9�9r�L�R1�RI�C�4_LT��]�L�W���=�V��V�qC6���������9�l�P�̋���D���E�bO_d���eK/d��7e1�Ç�m�Q������O�Wӣ��FȎ�T��X��0t��K���4�n��Lo�������l��X~"��Q��^�b��ba�B#�Oo��:'{����v}��m��[B�1�9�v��X ���&Z�J��T�v�q�)b��Ɓ$Nt�̖L�zi7�x,��b��bvW��v�|���t�������������pw�l�;2�+��0/����96p�
�j[��>��S�rR,W���<��	v��n�N�[��4�_Sxa3�R` ,l�y
..eN-
������r/-f�j�;�	5�&�t�|��v.�2��f��UJ�h�&o��\�|C���>6�����m�T��S����ò�a��m�����Ȅ�L���t�m)�yU��0XS[�t�\�
�}��x�����~$S�0���rS0W�Y��:��������{�(r�X쑦=��m�Dj�s7��� 2��͵�ރ�:[�W�1w�;&_ul���]T��	ZQ�A�@eo/��<"�V��7��p�L������eP�J����'R������OE��K �Z�U����앐	�����F9�_��~1���,�d����WS�� �(�Zc},ĐD@9�и�s@�y��w.�tb���!w^�1�;�6�����d����V(�� >"�.�"���}�섡AH�Vכ̜=�l���%�C���.m�KEJcw�˂��3L�ؚq*\���)j��]�h����Nt�$���X�F�{`���@�}�w�pp;js8��j��K��AI��ZصBddߐ�m�&��={�9?�[�y�F�nKS	�9�%8c�f��$�+u	|<Z�����r=�u�����u:���S�gj���i4�s��9��c_+i;_H��C���O��'x@ֵ���Pʏ���MZ�YB���7��ǷX�ך�Q����ұ��/�m�����	��N0v��v.Fi8w-{L�4֩wޗ�CA��o8���ݓ�6j^�v�MC���6�b�eY�O7)@}��M�Ǣ��K�� "@�A�[�h�����Rd.z�B�����(-���ǰ�����Dm����������aBG�,�!7��bE?F�����_��BZ����)��_��P'����s�g���$l"̓Y`�wA*�W}��2�5�x�(��/��[ܰ�A3�ٚǓ�P�U�0t4��o55T&@ ���a��}嚽�q��G|{�+؞�����QєA�z[�O���V4��R:A�� i�>q ���=T9���:���CѡS���F����,�@��=ۏ�� �*�
'"�wD��g;p��}w1�'F
������ E��,e���@��Q��o�w�1ES��a��i��գ��m�,���Z��'�j`�-��"�&�REi`��)F��Bh����j��\������&I�`r����"��+qQ!N��MLb����sw���Y%�(#�lU�X�� �Tw�����^��ŝ)��)�vz���}L�����85��L� Ma}5F��I�����]���l��������}���0Ho.��ĥ����$�v���S3g�}��ߕ�V��d�q����%�[�֡�%�>���� ��S�H� �W_zJ���HғS�P�/W:)XzĪ��x"
�
b���q��/*�W�?��-��-�#������U�@����So�^�\tPF6��R�ﯨW�겈�H�,��Z�S���R��{p�L�%]ً�P�D�����sǘT��Q� �(���sa�q�ш4�����+�ʎ�j�<5�R+D�r��d\�}����Y؍�V�s��%ъ�z���/�l��y$u�(>��'.Y2�(���G����B�i�<jе2n���r�V<���JS2�V���qı� |�-�p`7I7�:�\�����LzZ�%JB��;��u�b1��z*��@�������;�a�}��w�����n:�V�H�3�It��$`������z��f�?���@����_�s�VE(�{�x D�[���s&�d�Y\�����D�W��n�A9em�����dV"ϫT�se�� �����-ڠ�b�SEl"@Zh�9���Ҫ�R�Ν�Zga�6օE%�h<���:ςW}-��`��Lj�w�;�������-��Q�]�������6�+�I�A��4�c~�L�/+�<+$w�a&�r�Gs���D����-��)�2A�&�!�M}~����G�]E��L�X����%�|�z'��	�z0д,+e`�#wg묘�S���[no%�Q�3���]CQ�Ռ����ڜ��3jpNd�d"H�ڸ�D�L,�O
�Ѭ�D`��i)�՝��S�:�vld�"۫�[���Fk���,�uX��`8ᖑs̃�G5�m�Q��
;���h��sG��rX��NW��?�{���@�x��=Z�@8Ud��lW#�P����	o2�G�5�i���V��90����C3T�����Hě�H���0��KpѦ�M���e3���2�8vH������p�
��#���o�!��	�)�]�7&�����"��sy����c>;igL
I;���$��ԁ�&J\��K�%���|C�n0��|;6�=�nA����i8Myz�ꉠ����i��Z�_�U���!�:@M{ܮ�.2���Ɗ@-�/�>τ{�R����L/s��/I�B�G�&�9�ID�_;��B]լ"b�����Q�����x�­?U�jjtj��@J,�
�tﵳ-�
/cȱ?�T;��gC�n��R�fهM�H�������6Å\V��=^r�P��y�r�HRV&��i0��J�V;�5��
�tt�������}�ʄfձ���~�ݐ�õ�56����ffKσ6����n_�0D���{o��r��c�X��@T�=�,���i1hҒ�C��x]%G���^��(*ũ��7/p,��<-^ �\xR$�;���f��PuTl���+�k@G��k��]tt�K�>&�����xW��;��T�@�n~�a:510���?-R�B��6�,`�+���6�e܊��R��o	w`g~�#��Y��9!�x��3d;��y���f8�aO�y5�&���l���O���;�:mˀv����է��5;��(Y��a ���<�kL�s�/��מ�V�Y%3<#�p���]�*�-0�����r?J鄍Y��#fH�?*�.��7��J�h�<V$$�|9� ܬ�vb��3��P�����Ǻ}�N��t�o���b�����0_!���PӤ�/�U3�$���i��LBB齏�@����*?�1%w4#L�[��!<�Q\��2��-���%�Ǎ��o=�ʊ5\n�̿�����+A;��?W�ɘ���N�h��2����5?8�l�@��������ju&�/�Z,��w8oE�w?�?D�)��=��ky�2���  �b��KL�VW�'��W��CU1.7�"�h-�'�Y"+����4��Ξ����k��u|�J�kXI����KG0���m�K�?,9��p��K|5���/�;Z.u�{�g��%c�j@{h�O~/a^���i5�N��ԄeAZZk�b���<�[�ygvi 3��*԰�[�Ά�^���WE
������͒9��I��d(T�";
;��X��&�[sn����qO�'�{ ����[�"�S� ���=8P'�郒��#^U�M��UcK7�%�!LV����+�;�Ӱ)�&��Ř�IÓR��Lh��ޭ��p-D�f��o���g��=�E�B��nY���(�͚�j�@3�pWĞ����3UC������߯��pv��:��3�7];�oJ
d�1����ŧ�Ё	nl_��]���n��;&��Esv�xo�s�0VC�*d�Qr�)}����Ҏ>��W%S���X� °һ��wu��GR�6"h�T��ˮ��u����:��O�w+ښ|4�ôo$B� �ȄJLT�#
ʔ��g�;YCd#��up�F�lw��P�2g�nB��,�����N��>%P
�d��#H����;��"�h��xgŮ�d�c�0ITة싼�����?Y2$PU�)rK{Yx��>�՚�[@���2��JA�f�!��G����?1L���"Љ*^�}D��6[l^+l���%��H��k;\��I��#
BJ��=��.�,���z�]fc�o�`}�"`#�!p�+[a�ʔ�L���2>�k߻k1l44��v���k��a�'>Zxz���bO��Q�ǲpY�0�"9�9$4V�`��u��^��T1�IB�L-�	�ɣS�\���2a��)��#C��aA�^��/��>�����͑u�ל`�Y6��ѿ���ϤY�r�
ʬ����aG̱u�h��S���Hh~37O�d�#��y��pF*#�>J���y1�W�2-�:�l�A
ꂰA{IXBV���(���-m��,�A�']U����.�j�!*U�ȏkꌮ�������$[�L��`�8�����?�ۘ-�o����S�މ>/�A���W#�l��0���`K2I�\A��В�%�t���}��tg��g�pnR�g�n�K�Ԗ<a��K�5[��I߻�r�B�$���?���05��'hS��k���z�Ʉ�r�H���u��I z�.|=ƅ�� �[����7��������f��m��n_�n-Q�)�	�au�1��O�K�D��}�������^~�4j���x��S�Mj�ܺPO�3v�S�.fK��dC���E��?� K.(� ��J��x�1�G�����������7t�L��ݕ�?��k#ˆ��'Q�d�?�%�� �R�1G���2(��⋻�u�x�KN��O�����
�G���;u7D?��޻�0���}׺����N�� �}ͭEmb�g�R���C	��)�D�ʙ.q	�#LM
7p�. M"U�2�)}җ���k�aZj� �c(����e�����L���Y�!��K�Q��یcUъ��]�M����3Н}�}�n�V�#.���V���Ç�UW_Y���\{������v����>��9��ݛ27�6�p��.�@.8Җ�I�,N4msE�Ǉ�tG�]�ߊݭ�'�9���,r�~�I;���ȴ�9�v{fm�}�� k�@�)�=/'��V���-C(��ʏ���?���)������m����4�t��q<,ʻ�W�,�UZ�(�PEwI��U1
�Re�;�}�C���b �ZL��ߊM�Y�F9����D����������s���S� o��%��^���a����4ӧX�w�Qd�@s �~��lB�)�(��v��ݓ���6P ����X�5X��*�����p��K��*���2�hJ|s�"R�i��0��i
Lu��L�CX-��XVb�WSXQB��1��dL��61��r;&�iDl�p}-�o�|h!!K�F����C)�j��|�
|AE�ԡ�*Um΀�����}��`x�C�ʑ�T ?�ȳO�#����<^D�/{7#d���������BJ6�x�����|�j�O�5k�a5B�/�g14���"�#�b�g��+�����}N\;�,������̔
��>W׿�_���\Gv% bS�|r�]���J�2��m昽����!����#�Ҟm��XlxVHYEB    bf14     c60U�`�@������c���c�k�Ż�mBKf�Y�n��F���v
�&j��'����0�D�~<�|����	�&&i�OO�t���,�q`lQ5Dr���`;����+�e���ރ/�ضay��m�fQ�t=]���c�z��sqwF�n�MN�t���2�n�{�B��Da|j�@��-�Cn %-I-�x9���la	 k�{:�p�c�3��k�w6'7<��J�'��YVo�����6�X��ȏ��+�7fd�]�m�1C6)T���_Q��D�3��`1��Ro ���!rM�{v�&��ttZ���ą	V�Rf�@o�s	������<sN�!�l�(�^�[�W�ė@�ZaiA��o4�7��]�a �\�ٚ�d���!�(K�-#�)����+q)�a�|��,^��K��&s�j���|I��6�܎ �8�+�~ �Z�ж ͖�OL���ܩ����A�;=���t��r�6QQ��CB#��\@�R��'z23i�OκI�b<:�\|	spx|�R2;���)�Wm�d��C�Y���ߍX\�PD'=/��d�@y$'�$����������CH�f>=�8̨�� �8=բu�#���4��hl�S��7
/�T�a�_^fM=�]���E��\��F��G�V~�C�y%,#D)w�A1p���T����}_�Э�Xc�*��n]*"U ���a��Lz!iI��i&�n�'N���B!����g�����E����u�bַ��z#��^�4��F0�znR�����X{�Q6>!�l���n�Wk�?gp_8 ����E���.�e���a��G�I��NB��]��j�-�a:=�_�n5���v@p���Xj����L�G^:�*���+��$��E@	g}m���٥���}P<��#�,Yٿ�߰���A$p� r��3̮�K�a��~ �q��ʏ<`	�+̫��/ڼMW/%��������ɫ�s�|�/gB�ו�2FT���4�.f�/�0JT���a��#{��r[�W�p'v���C���� &6��0-𾔋��ўi0��[e����;ysК��f�����"���G���A/��i��$��R��Dq�����B�����].��n����Oؿ�Ɋ��*�������[���n�2_aj	|��3�0�J��+!�v��0z-�E*>��w
n ƾ@-����CB��0�l�m�����ޜ_�eL�q�&��7u<��V{ND�5۴
��&�\��|����&���"���x�"`q2�����8ّ�{���$��e{��Ӭ�m���4�7��t�
�y��x���0�C��`�E.ANf���8��h�x��t�d��ei��W��%<24�^�&+ʾ_���N�� ���`J�U�p)t�*�wK���v$��Ƅ�p���r�����?���E�GV�]'M�����U�6�'��Y���؂e���H�jVq�eؼ��Vbܟ}e��3ᓑ�O�Wm��4��W�����(�B��d�
��^M�����<Ҍ�E�<��V#�e�m�5�s쌜ڹ|�9*����\N�����gl�՗ZߤM)2��C��kGts	��[y��l�t�B�w�4��t�I���0�1�l��Rϗ 9թ&�8V�Q<뿔��[}&L0������y_##����F;92�&$82���3:S>2D�<��"Y��)4��DX�B�(:^�l[�e��2=-N�`ۿѕc1nn�Ϭ�uZ�%�A��=w`�|Gr�Id@Ĉ�� }%T�~��N���%�`���F�fkn��5`��O��㒩����׉��E�:�tl��J�2p�>�)=�\�6WM\� ��7�3)@2��vϾ�J�$4IQh��?�i쾵�;'e�b��R�*Β����uֈ#�z)B�ָ(J����D$}Cl�O�B y�y2L�)$׺��։c�0)PW=LZ��zKޣ�#G�GJ��[C��
�� jX�JZ���oQ�1�B��u����+.GǊ�D�}�~h��8�	CSV��o�_����$]K-��H�AYAI]00�%Y|�+�t�&�w�"/կ��e@����y��=^��������h����i5_�j��c� �~���}�)/mm�8�rE�m0�����z@�~BhN"�'�Z�&��|��[��o�!��"| ���KV��n\�zy�+Luu�WF�n@龠z�AFk�_�N:�T���C�QyO�x�8��j�ߧ[�$p�F���h�MjR�LiF�f>������J^�dg�(��b�!��wC���y�*r�%�L��z�����	�-�d��,M�}�"�7@Y
�<�FJ��:wu�m	3�w�h]�:eMU��D�"ϴL�/��I�Ln�wߡ/Y[)Sk�uh�Lz��2����h���qV` �@�e01�q��v�9�+k��7�<�H�rxL;��J0f%�\) a�?��<{�����Ϯ�������C7x�f;j�3z�iF��e޶@t�5��d��)&E.�i�>ڜp��_��M��۱-9�畽JD���&$�]�Ł�]I)a�j3ח����� �g�e�ӏJ�9[#��5M��K��{��B@p�6�)��6�x�J����&� S3�4z�1�?�?��ont�g-����2$���^5PnHuo)B����[K�ق�q+9Iv753b�1��H�lL䡋tB�zy hn6��b�K���S�a��6[���8xi���������2���L��S��QXօS-�h_�2e��wV
+a�%P�����3]�gXG���j��[+>��n�����a��<0(�at���n�o5���\��;a��)Q��`���A�͡�}W)��L�gs�i�m)��X���O3��]���︨m�-��8�i.(����n�`�m��m�q�f�ר|�e�σ��Ή�-U&櫖���r��4��Q1�����^�6I� �	���Z��&�����D̙��[��*���?F�>	� �U��R��M%�?��埉�R%=�ה	��`�;a�$P�n�������{�����{[� ��9������҂��
�i���1�| O�`8��