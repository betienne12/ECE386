XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!2��Б}����:�W�|ሖȑ}L�n�X�c�����S�V����N�In���/�!x<���;y/g��3"����I�h[�	�.xF�nS��00h� �1�4~��հ>�
q����D�ފ_�E'���#T}buLg�^g���{��k�mDx)�B�nnK]�o���s���o��v}��y��Ki�B$�,�b?ɲ!���_�MB�@�d��ײ�`��a�7��̉��\��`��X�u�F@�}��E�Q����jۭ ~���W	0�]��x�E̺��z��N�����K�,G���i�1���R5�]�Qܒ���'��-��ūF�ڄ��cc�=:�#� ���� ���+:���YF��`fJ&��%$��Z׀'����@�p�˶s�#���+^Q&����8�,�f�bG�?݂S�(����&[G�lx3�Y+"�\��*0U�JV2�
���+#��w���et�5._ٝ��ZW���9N<^��:�c^�K�w0�r"��/�-������{����l��L�u̐�Iy�PB�B"�da�yҿ�O�L!�X��X���q�t�L�A�L����R���%��ۓ΂�yk�C�x8�����8v(�$����o��c-rZ�FwL_^��������B���U;Ҥ�X%���2x�����C��j�ޑ��b�3�bf"ԣP�
;&ʺ���`�I���D,|����ƅF5�9\+��>�&àL~���Z���.i��ĝ*8��u���XlxVHYEB    33bd     c90;��W����1��t"�5��w��H	�_�������:z?����n�LjP�vY��,��Qs7��V�"��`��Gu�Y���K/*�`[^ƏẨ�\�glҜ�ύpDx�����HMY[ ���Ҍ��	D=�[�yc�v���f�w@��sˮ?s�e������ŧ�[�P�Z�Q/��DU�)�\�$�Nu��	��p�a�e	L�����F��f���tw�
ف��Ny}<�R��^�J�-�/J�K�+q��~eRaSe��yN���n�������Qu��>��uA�c�ⷉ/�(��Ƙ2��-ە���]K@�2<V�1�K��iJTY��q��	��VWU��b�3��:lz5?�*�@�%hCt���j������~����;ƎR��evI����6*�i�<������|B�2j�M�O�[��UHL_ʄ#6�����lRB�n���u����;�Á�n��\�!��M�7�#��ɧ��<��X�0�^�������I?�-��+#P/����$��ු��h%|��e9  !�����J���ɳ+m`B\M�=YH;�"jh౉H���O���\�A�M����`+��]_�"t��~�`����Z˛}I�D�pؐ�_'���>���l@���R%Ԇ+Rq��&��
�d�J4�Rɕ���Qrͧ�t���U���7��	�t�W���O 3qf��*ε������Yl�l�ނi)4�ٕ�1�O/bP��\i�_Spf�]��^v�7r܍��$�x�\B)x�|]�N��I{�́#��p��(oǇ��/��ه����O��N���6�q.��� �lL܄��������<L3pm�`F	ly=�C�J
!�Hp-�4�fU��P��U������H�h_^���8z�%�0�CD!��*�OPθQ�F7
�V��iQw���5:U�x���L4f;���h0�a��j��响�x��	Y_���k�;�^��񋧮�x��2/8��j�p�1\�P|�xqʥ�=7W����s���{r��Kҫ��O˵j�؀zi�b�!�EP]/��K�xx�M0�X�մWC���;km������f�!��+��m�00ꝁ�b7�r��Z_�q��c��
��Ѧs;�:
P[C�aI�5�$C��ï+�Rl�%�AO�S��u@E+f�;4����{G�w+چ퇆UB�YU�'�x?�	���Y����������Χqn�V��429=�VV'" T^ҁ+?��m�{0)O��V��)8�L��(^ ��Lf�xf�N�:P���K~�[ڬ�?�Wg�t�r�pD��a����a5�]�u�����.��.R��T>
��?y��ϩUG)ڂ�֙��>`4��-4?A}��m6�t�X�Vr2l�5蹮^��hN��#�r� /�kw���{V�D��khj�m��v�H�C��L'&�nU��� �(���dѡ�|�q���+)JΓ�D�lh��V:��A�e���X�[�Qc�1��{@����9QX�N/�l���.���i�"\�d�Q��}:����_��Xx�toA���QBv�7�b�<���	�H� ??Ȋ `��s�.g�3�������e�N
��DΏ���Y�jtJ�x��-�,=�Y��F���\عr��ǌ�'�����R��߱6�
���$�M9�b�}^_\�����F���T%�=2�
m���X��X�v:���נk#G#������R_ش�ˆS���g�V��4����f��&����	���%S�D��Z5̪��;�n�~���Щ�	.�:��rR���9��@Mm�ybg}�4(�rr�'�I��<��7��^���=Tf�~UU�f<���]Om�L�3�y>-<�J�JK�`h��x��qW������ID�:��r���!�c��>P�s�l�L{�0�]��%�ǲ���
�֯�����`%���u0��\��i+ֳ7���ֻ�/�R�;Z;Vtf!�ct�T�
������"͙ᠭ��^�A�Ih*�T��l�tUmG�0W��ַw���<��/�Q�>|u�0� $�ӫ�0����@��XH��m��<��]�dgQ����
L����=���Q��O-Mo,%Ҳ)�=���:`-O�1m�@���r[�x��ؔ�p{�`������01�$�&�/d���OTk�j`�u�K!���$���4����W��cr�T#I�������}�WS�.#.��k�$YS��� -�[�7�=1�JWbp�\釢:0S���	E�
P
��^{��A�,�v����VY�˪	K�Sv�3-�>�˲���W��kcs ��Y�<�(xS��/Ŗ?Eɡ�qc�v@~(�����S2Y{fqx��Ԡ�P�o����� v`���}��J>['�p.�μjB���S�1 ����U�H�fg����W�D\<�Y�߄� �����6K(~�[ؿC�R���ݫ�DY�e� �r|A�`�������*Y��|Rs�T���D�2��C��[�|�Ī�}	���k�b���� ��OR������l^1dNv�<5u�y�Ǧ�*�+=eVLBc��,?����P�x����ձo�"�9��	f�u	�%s�(t�-✗N�N�l�Y��m�1�5x� K�$�����}<B���n�{#1��{2���Ď��5'��r�*D}�%��`�K��'��U�2�$��<�2?�����ͤ������$Y^8:0��{چ*E �Պ|�n��^m��0�Dl\����Z�.�;%�Wl/qsq� Ex�ͅ��I�m���Rn�.�Tk�Q\�n���%kj��0�o��Nc}2�ĻQ�?�2ut��ֵIc�qY���?	�qB�ۨ�����I�UM����FJ����1X:��7���� �1y=0��t��H�:�{(Ħ?#nj ��9��a���[&��A��bm���z��P-��π�q|�Z���d̈��IB�U|j��Y�kb�%i��|�R�wX�gש���y��~�L�t��s�����j�v�E�s�������V9i�,�ʱ"巘�`�.U�4ּ`5��:��Y�Z]�[վ�tX��	���?�k�Ng�GΓ�."���t��������Fd��^�����Q��&0e��2�