XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S$��8���iΜ��q��S�#�ޡq{�a&*�\��캆�b@(�j���`[mR	�#��W��:�~1����П�x.җ��$X =M��bb�!׌��ݟ���1��(�m�fg�\���K��?BM�� ض0��љHؤ	!X�+t����X"1�����$�h��.#�n���6�lB/�!k�H应^I�i�6�Z C����c��Y	{�J+��~5q�M��h3ؿ��k9�������/� 5���~�}�D��]�e��dhp׶�# �7;Į�ˢ}�V� ��jG�=<X�J���ی�|�;�Q��'W��]��� 8�-���
O�h���TR����' d����4Q����U��3M#�"a��FB��Y���g�� {1oВ(�D��cN^�ve�*tK�ݪ�VքI^3d���G_'4�S������x�7Q�UeM��nɇߐ�YB��B��b�H�d~���F���k�v�)��W���֘'�b��F�Ge?��u�*Iq���,���n}t�=<ZǇ�=���ŀ�_��X��S�����뉦�(H�� �Ȼb0�4Xݺ�=�[a*w7�+�6�� -��!�]7�I{�Mu��P.r��6��n$��B�@���-S���ܯ����.����fIv�}�!m?�>7�� �HR�a%�ix�ȑ�[���'��2B��C���N��&3Ћ�x
���3�[���RHʆ/�q��P�v� i_�4�(�˅ˑ� ��XlxVHYEB    aa31    1e40h����+H`�-:+t����,{�M�?�
m��W�NsD�-@��ў	��QQ�hD`2�p�E�x_3�LD�U��s_�~^y��z"HD�J�h́�ݽ<���;v�ci������crq��i���b��=�d��\x�v`~�=uZZ�^�r��q .7��-`��k���Ej�!�I��W�q���}��	WU�*��9[X��L�RrA�u`3Q��)-9�m�Ve�e6Z�;A&����tF�!���Ή%�|�����,��Z(��8��v1Mיk���٭����W���!|����}�ˆ� 'U��4ݯ�U�sS$]��;�$Ѥ���:g�Tg,�g혊����E�-t�a{.�r��2"�z�W�	c��A:w#m�-��ި^~��8fo[�۪�Er
ň��=9,���&BXe�m@n��2CC��Y�&��N���as"V���홍�<�p�{��͝ ��@��wrp�K}l�N�wSF�U�\WK�r�u�.���Ӡ��O��� �W��Ś���E{�v#��~�D+^�^��K�cɓ> �ѽ�O�v3ʥ�=����K�$�8�����>&���BU"�޹J.U��>���L�uLw2����oGo��e��˽n����_�ᗦ���h�͸��h�B�A@to2�%�?���l��@����v�;�:�+S.���0�?���+nO�����v2��:��gڀ�mp�)�x�Ƞm����J���^�VDDu=��(�| =t2��Gߋ�`�z����p뮼���6�u��c��t�e�%�W+rq�<� ��R�7�HB�Iq(�Yݐ�G�N��&~�yg_�P	�}�m�F���%�|+8�7ϕGG]T}�!��Oڅ�h,��GWۺ
5T����G
��"ނ�j�X+��׳=�/�� �7*����-xi��Sh���8"]?�K�j�͐�z&=7%֘�XY��ɞ�QH`�-�0�x���)үI�#:��"�hr�g�85�8�f%{�e
6W��E/�(�d-GYJ���^����Lɴ$��]6�����D"᫷��^'�= Bo@�O�v���U�s��fk���\UcA��� S&9W���{ͤT�)�
E��,0�7�n/�% �EÈ܄u�"t��#t�w�vˬ!��\�u�;�B�����_Ҕͽ֐	<����%�g&(fc����ƣ ��&|�sp/`�%p��0�������\"��jS��+��Y�}��}�F2��1EO���ި�����mgi�����u������@]lI�(�"�hw�2+F/���#XIܜ�wF|��򘳋ĥ#�O�0��@*QK��ZVA���3.�yrB������]� ���$*䟅�E�!�nt�/���O<"[k���䅦��F�c&;�y�_vda!���k`en^�4���bd(�8#;Lmp���CK�J��5&*"��'s�v{v߉��"0����~��1�'���~�������WԌv����G
/�]�
�!��%�M��*�)�7�f��.)*d�X5��Y���ȰZ̸ܾ΄��3�Z!XT�Q��箠����m� 4?���^=@<b�QԎ2t������j���Q
���h������jͭ������\*q�r+�,���\���lT2�+b7�av��.r�%��%;v��W�:�W�P�,�PP��ZJ tCS��1�� }�þ8���j�KtK�= :Hp���0dTN�"�-6����zi��u2i�9��fsed���s���*D���d�)�'�1y"�T�J=�L~��z��������_#��EO��U�C_�x�v��#��s7�U܍��TE{�܍M�+��>�7�D�tҹ�W;aXz�4o�a�## n���:�q&l8}����;|hM��b7~��53� ��Wo*�T�,�����\&��<wX���&ކ���_��o�<H�r�����Ld�:8����Q�n&�	z1'�8ޫ^�4�	�RmaƸ��vZ��yڡ�&]�,8-�xJ�J�0��	B��sl:�s�TZL����@'��Rhfv�d�77`9��~E��z�ʝؐj��5W����紊�"�pʩY#ZP�	HT��}�V:H��.�v#@)0�S\���w�/�iG�{ oM��?$�iL��_�y����jk���v��U��A��h_�ݛ���3�>�vj�e�*-�VM�%�Z��74gL���xQ�N��E�>�S��]��@��'V���Z)~+��,��d�Q��Byf�f�Pe5�BPK?���$�����lO��p�E�0_�	��$P��GB��jT�����T$=�o̵AU�<��^������}pmA�t��(|�'�q�����F��n�!�#f�|ZzM���6���4�`ǰ���t�z�m�� T�9dDLyQ3 'Mw�-�u����U�g�g<�]��J�/f�ow����I��čo�g�H`���wV�0A�?�f��p{C��/���zՆO$�)�2e�ޏA�ť�H��5T!�"�naq�0u�8�eS�4D��a�,O�/�e�jL�|��7Ib"�^����`�l�@��c��:�����q�q��a�^n-"�B�I����={�60�R�ƹ��U#�2j�5'�f�Z�~�yl)v�Up� WX�7QK	��4�32���Uw8�e�
����W�5u��*�#_ByU�����8K|�D��*�M��R�k��Q�Y�#R��O%�Wb���!����&��L�ڛC�#���/�pD��q�c�0��^�(�ۚ((���X�#��]dPyP	�%�g
��o�7z2JN��6.XᇆqpυKX�j!{��_,%J���GU�mH�R�]�%_j�}*9�G��OYY"��*ix`�i ���j䪩�r��nZf��������	�U�,�1B1��&�%|-�%F�^�I�<�I�"GPl*�6�R˗)`��-��a?����o5&ѳ��(��>��U-�*�k�#��izw��(�h��v��H9��9�1�,�s����!���R@p^6����Pf����570x"��|̦fj�$��{N�9�̨�1��k_{�.dSB���Ҫ�!v	�%��#���B��#����N~;��":�QS����W�f�p��c�����u���k�r������KK��}%a�|� ��T��g���N;Z�Q3�Μl�"1�T����s�椹��ɡ��ㇳ�Q�m�C �a��>W����ܢ���T���%���9�3��jz0$Bu���f��0����:ի��x��+u�+�4�0�j�?Q̝ܦf�����Z�L=���p/	�I���u�L��;�J�Es����\\L5���p'
{��lq�˖5��'U�O^&�/	�)�Oy������D~?+��n|hYU\1������%;Yr�������l���<�і�K�A��O������弎@��V��Y�|�����	�7�|�8�y/�;�a��L9�Wy�γ!碞J���
�Dbg�)y�;�B�0pz~ 6kO�������8�*�H!]��D�U9��l�v(��7t�v�}2JH"�l��qbߵd�$���	�i�F���ęa�x�g��Q�xV�Ǡ��� �g���=x+4|/;���d�M����('s�w�km�R�h�[�Q��C�%J֍ex��<�
�/Y�,A,�����h�/�������^���Ӂg�իh�>��JGqX�l�{�<�	�����-j�\��6����g�~���M�`���=Z�C�Z|ϖ�9[(U*�_x6�R�cX��v�[M:[���'�i�S��H�Ta1���0������z+��d�L<*��	��(+V�խ:�Wjuq��˄ރ�}|�P�&��df�h:���������	�;�cD+�;٤甴1���$�H2�T�E*s)՚�mT�W��������{�R�dRk��W��<�E���|G��CS	�c܌�j?)M�1i��C�sW	:�T����ou�3^e��Q�g��rWvR����";�- )t��~9��������Aq2��M�u�C��g�#��۳Rk��r{�tZœ�O7s���E=e��F�cƂi�w����_���B����t��t
Z�+�Cw)�Ғ�,)%V��,e�-�x�x�r�W�C�R�#Ex�g����_r5�7Z��a�Z8�fD�ύ�5�-hX�гFx�=N?�{'�~[���{G��\}	j�Y.S?��q-ĕ�WnJnp��C �m�p!%4�Z%w�����S a�ckm�Rt�Fg��1YR�Ԇ��h!ƃ�?�K��]ث���?er�W{%�b�8q3�5&�՞�F�ڞ(|�O�c�.%�����H�kɋ�� 1�c����n�Kʖ��s6R�/a1Dt��W������ĻPa��U������-��9�Q=���@�T��K�G���#�Ӯz�T/r��lx�O��a:�(�o�������l�L�e�x34f��*����9�#9�=4	8��>EtX�]��̆~X��*�#�K��U}$D�tґ@@������GKIF�h�ɳ[(�a΀FA�kD���qmK�����f�[d'��(�[���K ���+l\J.��g�]uls�(Ê�����9I� ��П������^ ��$�MF'�1z�t�n�G�L�V��TP�̉�8C�1���@�1(���SW�G��I�W�\&��x�o\�.��S�3GH��F��A���/�w�2�[10�!I�i��-�W�+�&�_�^M�Ҟ�+�w��3XZs�\r��}s$�0���*\�w����r����K����T��d���J��t�u�Թ�l�ZL�V�Z夔�-Ů�����h����Z?�t�a3p�|�*̽���U�=�nb�e^���`ĳ�G +����o�]�T�޸�K&�Ŗ���#�2{�z�kV'&��T���T}�Zvg��HR������#��˻�А�ew�h�p�tgׯ���A��"��r�b2����#ƺܑ�G>�ݨK&��z���m���Y(MF����"�#wfs�0Kee-Y�h�v���N��0�d`�"�ʄ�T�J�(%��a���� E��]��l� ��/�c�7g`�u\N��',j9�
~���^�Y�F.�����8�~B��X{*�=ů�����䚎�5��D����}�,�P�]`r�2U�n��H��h>̳2]`�����S��D�9&���w Y'*�B{�h�U�r]
�b�YE7SAAwR.�{Ā��	��:�P�,}ĵ�xbu��t�G�h<.��/k�4+;�WPyFsCU���獢�� ��������75IH��dp�MuN��M-�K�	��ZG&��A��B3�2��o�#DKñJ������!��i��8������I�Hg�e���6j<bن$�|��ѹO��8U3/���"9�y� /���>�L/͐i�ĥ׮Td����U��״��N�{@��׊���ُ�ŧhb��_��_1-�#�v�lT��7N��%�V|���zc��=���np�s�y�$(tȒ?�6 K$��U	t�*����ư�� �F��%U	7��rx�����X�����Ɂ���
f�Lh�J֑�mH��Xޒ�3���%���+2&VA�}��B�K�q@43$�MYFy���ܑ��蓧f�47<��ݧ�]���=��:����&!�$�}7~�q���+sz�x�*n��#˦�P+Id`P��KWV�j����>���//}�ҹ�
��霑.�U[���-ˠg��V��+sS��@� �^wR�W�hl��$pph�M����x�+����0u%-���-�Y�,��}������/?jݛ�8�N����+�ulle1�4��"&9��7�:�q���9��4d;�!�� a&�_R�h:�P�3�W�D4ݮ[��U�>C0���V�R淋ϒ�B`]K����)�.��k���Y�љ\1�F�ѻ���8� ĬBjM��e�B��nͷ$��j��ʁL�m7K��
�l�������w$�q^�Ӻ�|�M�c���D'X+�h��!���l6�>w�u����{���S�p@l!�FR���3Q[�2�7�4��9o����!3�H�q%5h��W�5/��2�ލ�����g��+G"����ʛ�p	���N]
�,/��f�Є{7�T���ݷV^�ё3�%o7�k���i��"�\U"w G[�+g�ٓ�)��4�����Lvh��%$ˮ��i�#4qTq�U�������͑��wE���X���X5��Y�l�p�{{yZ��zz{���Üq�����X"Wi����$�j��Q�n�p��R�������y�X˲�k�����[��6���I�+P�p��+��#�t��>}M���(���rol��7�������?�@e�Z�+�F�("
;��F���I��V��o]ǝWl����U�j�q��j=�r�T�=�W�Uz7��lόt.��!�yNB�$@����,W^�s�b������_�O+�[y���So��q�l�iW�$�}��Ix�Z���C؃_7t�/�N�ZEb��l	����4�5:)^��&�Qb�S�s�k�BԈ�,���,�=〵O� (nK�����p�F���}������*SX�����MC�5�ԵD��_�/T���#/0�ԃ[�@�ZUpԌ�^�	Ζ��Aa�=��3��+�tzB�RTOJ�ɏ�_��R��vnh������Gw��S}�r z�ޜwh�#-�g6ih/	JJ�9��ʉW�B�f�A*2�޹�����3�r�qCޭ�*��˹�8b�L�xX�^,O����h$G�?b��g�&�I���1|Oe���oH1�FZ����|w��Vŕf����B�.L��rο�ii�����<�
��B\�m��HG��1?����D�F������T�2�7�R�m��_�NХp��FT��b]�gI�n�&Kα�FGii����6}G��OCϖ`7(�ٔ
����ZEK�[���Y�(L�z�����
y@^�A
r�l����w�[_�a����O��X�B��(�(�)�:O���Hz�abo��^S��_2Kl8��OɊ�T�R�z^���ĥv
��G�"~���R�;��8L 㮦�;�&e�����Ǻ%
1Ǥ�g49��bAAL�w�=�90�1���:���׼d���*y3���D���[̣r]F���=�HU�m��rv[{�#�ER֝�~�$e�B��I���B8��v�V���d_��x�W�H�-�q9��S�B3����YO��~t�fb�y�Nc�ֆ����� �N���2}���J	�E�`���;�NujK���&-��3��(��P�(�}ey��4hV��%407��HP	c�ꛜ�n�	�ޟ#FL�K�����.�~�e�Nf�P�y#�JiS�SE�L���R/��Z'�fI�	}�\^�Ư��Oȇ���M�ҍi�#�	&ܐ��ϻ�ĀM��.{Kb����8��:�Z^t�b���'�rپ�����nAř�U�vqӛ�h�H]�W����'�XH��S��n�w�!��Î�0�