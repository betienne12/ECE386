XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������>���Ǽ���`=^|�ss� ��lY�W�����o�	�l��|̆"�،���ʻ�c���ei�3 <8�,�#n��rU�)Ƣ
���{�g���L5�]w�X&��Fڇx��|������v/���� �b���سed�N�w��x�(ߍ�ㅢ��Ú.A�f�7̈́�[�����`J�
ў����]@g��٦��@Ed�+�@�i���X�롗e�<�Pw�\J�`h�ph�X?�iw)����?z��?Q�w���Zn�&�}�����FN-�,�e~<����'R�x�t��Yr��޿[Ϥ���\�~�����3�
��� �3�jT.��h�'�j�x� O9@�c���]PrΔ��f�;R���.�Ι���s��
x��,���C�v搃�����"�T�9�(��k��Rꤋ�DT>�t:�0>�o��?�2�0�7��Ehx�n���!"���6���$�� *�!
A}�|�����j�W��R�t�ǭ�J���Y��=�B�G�f����bQcIu�v�OkT)����P�	�&ݼQ��M:����m�щ��d�7��}�=2w��)62�����k'{S�o��nkm��A��)w�%(��^?��B���x�G\�tx�(^��f�o�M''�j�9����hoQ�*b,w/ �1��\��*�KV���e�K�5�yY����Lr�����:{<�X�<�OM��*�W�^"�nXX�S�����XlxVHYEB    2e55     b00�OHK�����8~yt�x��T�kϔ���*�C�"г�L�6�7�����c{n���9_��w.�0�p��D3īT�'���Dj� ���,�>���!�dbWo�itӊ5����T���2'Xd%ɬ���c�(@��,c��o��J�N��i�Pч㉥��[��߄�fp�G��e���͵�!c6?�.�!$&$+��W;��^1��>�/i��QT�ջݛ�'�­y��S�k�sT8&b�X��5�����X�*J�&�c�m�7��C���&�F�2p�ޥ)igӷ���]G�'�ݐj�ʜi�o�qIt;��Z�STnU=���=D�^���"�I)�L��i��#�����Y������T��1�V$i�Ȧt�(�}��Ϊ&EC��B'(}����Iya�s�M�潢�ecDv���
+�N�:���KB˾<��.}2����J �s��Zeν�M�" A�vW�5d?�B *A@X �%{�\�./�@��*��Z�.[�8m'��m�.���x���
�jR(�QM|T� ��o}Q!M���:&��mYeL*��9,�0U���w���) gQ�w���w��=�`����_��6IXPc�\h��G1��+#�
�Mb��Ѿ^���U�Y�����rU�H׸����Jn��w`׻溛ܐf
�G8����o�:�Dޭ�]&3�!s]s��Z��u���wu����|C]�^/*�q�bsg��TVw�"����ܿ�0ⰻ��7m����5��� �9���$��IQ
�ae�������*����@���i%V?e<�SF@+ۙ�ЁT�#Tm�����E:LBA�x��҇����i���,�֦��#g�}G?��2�5u#�&��@�xЎ+^�jf)�f�cm�"�n�p/
�fjpeM���Ś��BI���$��;ϱώ��q���#E�J%;�C�q'�M۷�0Q��G+�-��!k��� w#02�5��Xz��Vl��!���%��#�ZC�r�O$ц�����s����A���jU�F�n����>�������[:V�^d�ńp^^�`_:�����W�Z:����v��3D�k@����U�W�ʴ����y�� �'@:���0f*���#�Z4?�m
�/d*���?A�r��C������e"�L�����a�_W�N7�W���`�Rc�����O���>Ҧi��L��''������+��eB�� ��x0a���К�T�87�ՎG������1�S@�����:���pO���Q�0I%��� ���Ǎ������g���⏣��x/x�����%^���-�^�K;�ȱ��h��Q�|��#K�"�#I���I���QHm��m+��y���7�Г����
R�[�8��?�g[	��0��`�\#គx}�&J;����5��C#ǲl�y�W*v��V�[�G�&���3Yˑ��Mjֆ ]�>'�E��ͱF�)�(�.��t�G]#=�Bt� v_�<���	�F��7�Z܆����*oܕ�W)\�$�\_�)i>�����'�<_^�������Y{���ζ���'-��o=_�����:��7ʶN>�p4�������mh$Od@��W������IC]m��^eHx�1�"��7y3l ���0��/g�ɀ)=���&{�6�{�s�`X��1iEV[�����g���s���j�IB���# ��fgq����B��O�nB�ջ���n��_á�G�:���}���e�����+�gw�S�"��pJ8{��y�c>fW����;C�Ea�mqI��K~�����С�0��1�
��F��Җ��WF���ca)sQ��|G��rS�̵+/G�|��=��]�/�m�U	���Z,�j=
�m?�3�V�Zn`��v`&���pȬ%L�|�R Ksd
ު�z��Fa�ŷ*�-���u�@w�c��r&#����9��׾�_�V�#�.,)H�Q�`kKgx��t��H������l�;��`!u��i���Wh���I
C��O����ï�0���d�+�S+�SJ����ڎp�tzh,q!$�./��?����Vg�����U������fT#1Y��;�Я��v�3)20y����X��X���#7�~Y�S� �	�
^�����n���L��b�j�U����(C��{��Ӧ�W�NI�3"�|�*D���������Z�̊=���75���l�@���d�
N�'��J�K�.����E��v��(}��u���d��.p��`C��z q�d]���+ZvڗU�bjUr���(_l�D���Q�)p�GO)�^�/oQ�&�`���"LVT������O�(���V���#����t;����gN˶&%���r4�b�z�s�^WG�\L�u��g�é��D�:�ў��=f�7.��o�a4��z���h�'�h�[��8��(U
�U�Cfp;p���
b�����$o�3�B],�˃� t}�S�}ɖ0Z���"8����r�-���-?��e����+�6k $��2��e�j�3��=����U0@�5�]�Dn�*w=��R�I�n��87^�٭ɷ���ם(��(����$�_�sx��c�C����svŒ�ɼ��Vv��nrG�8aa3}��L���Kt�QH�4]3y7\�G�׉��ƈi��w�_~A�b{��,�*�w7krԝ�§��MI�-��]$��G���aP�Γ�7�����5emB�Wp