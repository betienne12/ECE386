XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u9�*2�����\����ƫhg[T5&�j�=��r���z4 �N�J8IR"�!�FR��RA�ȿM����\!#�Fw�?m�I������Z��t=��iU�ZY��ԤH���3�7Q���~����`�)���
S���DoN�̫1¸�-�Pٚ2z@/%V��bԾӠ&�Da֦��(�E�d����g�>�"��h���5*�/��E,O2��u|��|�0�/<�CA-+ͩ�.C�v�
q���:��~G�p+.u�l�C�j(*:׺��@<އ@�ajR�>C��!N�V��ex6ϵ�]ʭ�N�]���k��\;h�]���yp�>�^�r�����]�c'�6k�b��Hw���x���TZu}.���-e�Նfߍ��\ui,1�.��0۽�Z>HԊ�5غMp�����l��4ȩ�?�|���4�ec�
^��jL�7����0n���M+�b��ݛ\]�z$e	���%Y����!6��v�1�{�"��-K))�u�I�$\�t�|EJf�"��s�$���ސ��87,Og(�WF0���_������{��:��\��tc�7 ��WRs�͢��~��Ѐ?U�	�^�=�0U;rXμ�&~������[!������\Ló�Ѷ��0s?���._|��z�m�ܞX��;��{�!�����P�6�ؠ���L�@zTJx�)�y�m�J�_L��~W�!|3���o�XM�Nr~"�XlxVHYEB    aa52    13d0���عM:_kqˏ^��s�P����A����
\�x�<t�+��~�2J*�r�������sB�YӐ�A�ҟ޼�j]�1� 	1���uΊ�k�ic�*w7hYU� \l��������>9�]��X �d�$�)`��=[(�R����1Q+<�4�
Wم~�N��l����|�o
{#��@�e�0Π�[���H5�@�*�+J�9FV!�c;Q�=3�����A�|.���m�R���/�����$nb���/�osx��R/��--����Ņ/W��8�e=�,�o�h�3X�0T�Q.D'�r���X���!!7�Fg�6T�p �M6�u{#�	�T�x����:9���k瘼ըTO?V������I(�_����P���'�ѻ4_�����)54��8��҉�p�Z�?���*yΚ�2\�
c���%���!����	�l)� e��E�l�k�D�P��mpE�?�Ԝ%l��R}�_ew�:i7��(�l�+���B�9X(%>s"E;���L�y(���E"E@�B�W�s��o0��0lV�VS�n�DZ�N�E�s�1x�}{K���Um�-K/jI��q���}�a5����0��`���Y�� �kloJd&
,=z�t+��ו����� �ڞy����_�8}��?�UM����kL�Z����)V/�Q���H��qՙ�В"Pى�\�����J�Ja�u�J�!J�Vg�N�[̬w��ŗ�9�(��V+�&�u6�7������Ĝ��@"
u���~�� ���-�M�E��1u���Sh�g���������i��p����{f\��o�m����B�+���v�0Am<O	L<]�DA@�2U�I�!i��$���MX|W��B��i�$§	+ #j�\4!�r+ ���0���`\�� �5����P2~!�]j/���<�̉���-��F`��C�`�\�of �B����22	�t��<U4����9Y���)~�T;	o=x���FG�u���x���U��V��*̷#���s�3?!�?�5��fu?��ߜX9�u�"W�\.|E��?N�=��:��~�D!(�x$���R&{��i�M�p�V5j���a�h��@�W���1Ԝ���ˈüMHfV���顩�5/7h��p2�h����u:�B���갖���_?�F=����3���!F�b��@^�H����`���,GT�2^ѻ<]�_��E�t�Wr�(�D$vfAf���
t���a����P�]H�EӠ��iGW/W9��wy�U|g���|��n��Hw��_���~Cq�Ә��
7����f\�mi���X �SO��!�8�1t�b˻$�&��C|
�E�����q��kvԕa̾c/t� �$>A��y��(�0HfQ�
����_�%���/��4/\h�sλ��=@\�Վ4�b�E|)�sX���U}xb}��+�i8Y�돊�7!��b�YJ���q�W��jVQ�`<!kė��@�C��9E4�$�=_|`��8�ޭ��,����7��`�A�k�1�<���ҖR�iM��Å�[ sʤ�d�oIY9��ՠmp�s��#+���~�{Z�ÿ=T�dt�$�(�����I����ʧ��0wE1��t�{�L KvP���-����J7�j��D�������]zl}��s�Ɓ��̘�&C1�g|��ݛVe \C�U���i�����ל�JB���W3�z���1y�bʸ>ކx�s�.��8iZf��+<0�����!��5�r�vT�A\������4�[N�"��I/�*]ô���O@dꡅ�~0&���uǣ�im`��*i��t��{���A�ˀ����k��1�O��ZY�JQ`��29N������UI� pID�&�,����+b���M�of?F-"sƓ#:5�'p�f���ru�'�&����gn�/:SIv�u�j�i�/�=���<���*���Q�J�}Rk[`+M�%g�ɫv�G��m�5Ց~闱��|�u�X$-����*��A��?����͸����xg��Ě`�TMW:@�g�p]~Z�X�ʴM�����ʨQ���ԕs4�!��%�kݴz����m���\˯O"����(7�#`�h�F�8����@s};�:?���9��E�����O�le�$������`��W1XH)I�Q��2���.� )S��$�+���)qk;	.g��#[����;�`��r_��&7y <�4]�O�fC�λ���nN�!�s��[c��F����Ϥk�(�^��Ė�_�k-Ć.m��� � �
Vl��@��*�������a�U��.�xEF��¹�>?\-��6��ک̈́1���i�WÕ��(�h�-�E�"�P�,���-�����f��\a:��~.w%�Х�T���9zbl����6���y����J
��{j	��q �kxO����&�	g�kv7�)�#�x���z�� }�q+�F�Z#��F묾��h��<Y��c�H-q��t8�L&R��ܝ�U��:���u���u^��2�m����b ��Z �a�n2pF�jm��9��pg�=8B4�q'��;kLDfj~&�������2f��F�b���ʍ�F�d����	�TRA�1�	K�:]R��8���ŭ������ ��U1�q�U�����l�}_�+3�t =Pe��T���~�x��N\;�
�}�	�/�弒���t;�����ƐCsY�SH�'*��,L���&�uK�ST�;ͳ�_�~	͝�wg;��8-�'�?,��,r��z�҈b��Z�Z�}��:�6X�x�8��f����b�i,�����d�wOh��\�AՀ]b.�gh@N�@bPw��,p�(��z[r��c[4�̱"y Ъ����¼�$�!^�кq��.a2�c�ٷ6ٙ����L$Wﮂ���O�C�%��߆h�e�R��ｲmTE	�ݼ��|?�H<F�ok=�<H���ժ��n��Mt������ �T���u�Ai~��_�G� �fhE����0[֮���a�NA�:�Ju�����p�����G�/���Tѣ���C	��`!8mNr|�)�ntM��j�{����ӻ �b�� ��c,mr�o8w��
-]��D/��h���^�sd8����o(���5�G񈓭q���)�����,}�sm*�h�����&���"��\''}��
X9��r/�C��AYd
g�ou+���;t�����8��i��c��#�h����U`�Wa_���<���������F�ꮪ��}���7��$�tq|L��&I�c#Aj�Wv�f�m�aU3Li�����8��o(H�+j�"�P	6��������+-Pϊd:Z�C�){@bw25I�ݩ�����_AF�h�C
mQw�aQ�[s�c�\��}�x��ŝ�ulzi�%C��	ww�'�fcRZ:���>��oϵ������0���봯��I. ~�#�\th�N��i-07j����Q�eOˣ�U�����o��~=X�;\V���S8e�$���#ZKV�iԢ���5P��pܺصc����Ѧ�p�<QC$��T��$$���an���7K��o�Oby}˷ؕ=�c	)"��A]��+�U�Ȩy���0{�J���E`�73B����M�gR����;�
�Q�Y�R�/��шS8�7q �����x�H�b��.�l�<E@�Y1r�v�s�R������.���]�[n���k����
�H��ѯPު�X� L���%Ox���}���n�c څ�M�F�~t��d���em{�lo�o�B`��$$�ȶp,����_�#K�,4�@Ϛ��6`'�'���9����7sh�Է4��<A ٪��!��ML�Pj{�M���,��
#:�ɃRY.�{�w�U؁��2-��L�z�A[~�M�* ?opP�ܦ-���3"-�疰-��-�֘�\ۣ�
����C^��Df[�11�U�|y�_Ƿ
�X���8���t�;*��?{��	���=loP�9�˴1����8���=F���$����I+g��'��q�pR^�i��?�o�M��q絋�z��7���S�y�z.v�����p��Tc=LUG�5[�6�A����K#
��.t5�o��$5mH�
4(�5�����2n�QNO�8�2�bP�ѲF�m�l)�R2-������.�>�hE�[/?�6�,�g��y-�l�l*���z*�ȮM���v\�YoN�%YǪrYG����ݓ3��w=`VW	��n�~����_|��U�z�U�{����a��N�]��]���t�1U,vLu��Zx��9��Z�k=S�$�A�`z
�_T������X�m��r֚�W��7_uKET���I*T�֏��D�Kc��\B�"�=p���T���*�//��J���/ΪR��v_uN�՝�2dz`[��%�Ř��J|.�/"k�5�f�\ �Nf�;;��6�����G3�X��M��o�l#Q-Hd���d�<�4���o_琀��nz�7J{���%gr�����R���E��@�!wG�E�iyև9����'s0�x-�������=p���7Ã:N�5e�T�!�5*,qmWvRAT&#0���4��9�y7nFٟ�<�<*-$�E�fp$b��v��M�jԝ�U>�b��8	�� ���e�d�������t�h�N��x������c:f���E �K���n�K�
�xBAar���7{x٭ZD-W�E
���ׄ��d�CW�fQ�.h���,\8@�Jw5���~>�`�`����ѫVx�}��=[����l��)����/�Z=�@s�#�3� �v�ِWp4YN ,���S]~ˇ�������������z�<�������>�}������U���=��c�bM�'b�J��^m��	n`��D�I��0���J�g