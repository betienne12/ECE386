XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B��hb0r�����B�&!B��o�H�$�aVň��������B�M�20fK$���k�1B ��M������+��߀�ʶ�"�p�O�w�������_��6h��hq�����Ic�0ҜF���� �9"J�1ڬ�7�#�-�*�r�c�v�k-Y��^���E�LJ����L�R�Y�H�z�|�G�k���	n�+2Ծ��}�v[�{�V`���@)`Q�����&N?����\xV#�UDXB��d^`G�ky��f56���M�h\�P,�^�Z3�&�|O�'`%F��m*��|��%m*���Z�1^����uM@@��X@�T�RT�"����[�K�{�㉖_¶�?a�<���.�)�H�_�8{Y���cȟ�Tp����̌03jd&G���&E����t�4@������7�l�[�3wth�eW,M���jJ�V�h�t�AE��ͥ�*���Cc~��� h���8fI���U#e��ꉝ�&[���+�u��+�\󣃣,�[_Z������]V=/��M�3͒h�Cr����\�ri�`�&N1�����B�Q�ƄX�{mv������b1#^{R��y4��9��so��\IrA����
�M�rbn���?E���!����-Q��(��7�'_~�<��=h���!}g��M��*�6��0)�X:�[-���&���P-�˱2��&�=��˹��^��	X-O�*�`�/�(,'T_wU!�ʖk�Z��XlxVHYEB    56d2    12a0ϕ�d&e����7Ĕ[��:C��e�M��U���K��QO6Y�Sk�Y���|޶P�{�nTz0vq���|Hp���rr8X1�Ń�|��k�^ʘp)h��7Y�3}���GH�&q��YoIll7�gg�$v{�񧕏�QL�@���(x������eJ�8���y*�JI����ۛ�AΊ���]@ٲ�~��=y�D�)�1Y��%D���Ԝ;��V(h���k��ϥi*�l��RG�`FJ7�В����:2\���f���a�@�^3�^i|
e>6�f0�w���Y/@U*4��{�}�{��8\�!&!0���ٻ�O~�y�QG{�0T�N�0�/�)�R�IZ��qƸ����q7S4J/���L�y6?t���I��A�"i�Κ]3�E����y s/�/;�xfp�'7Z!+G>w���OqԻ�1��tPjxx�Ϗyi�U��$*�Ÿ�\4#�U�)�6+��k����`6��3`D��(&	;+���+��ajr���tm;+��|/��<���;a7w��(ZDp�gjW�\�Tpr�����~�G�q��L��Gd_;���ʑ�_�9Q��	t��!�e�{��ᖖ�_&\e�D��M��"�+�P�Ǖ�ɔk�����w�6��s�W|X7@F��%9$M��>N�*�z}�L��Acv�`�r�Мn�����K�,���Jjl�"�2a%��R���Ɏgͧ�-��ع"&~~�N3w�%�C_�r޻��
�0��K�r��G[�ƭt�ojQ���g�p���VX�=ze��� ��������>Ctж#R\�[	��ګbf5��'[0!"���$�k�Ά�,�K���Z)��k�-W�Ә^��`p�����8u�atɮ��_�,0yDv����&���h���f�Hnga�v�����2�������ox�M(�k	Ա�L�(�^̈#c���H:�gٗ��6K^�_(��	�r��Zs�1
�E��������V��b]+ơ��*�������|W��qD��W��@�K��a�y���"��ϋ�?Y�M�J6 (?\㫰�oƶeᨶ(=^�BY��BH��}mB�=��Qp��f�(�4O�r�$�r��t�%��#FL�v�� c�k��x�����ixC;�
F���%;8[R��z�E/_j�l]p��	�`o{��$Q#����XH��;w�%��Ԅ�H�Ə3�j�9�fRf�d�RY��J��J���'RL�T�j�)�4R���*ڴ�yd�4?u�$�6�G���z �^�A�:���:M(�$�i+�)S���-}���j'�k��&a�J�R%����. ن{Y����WT�#~�;��f�̊W��S�@T�E���9����zpY�J��]k	�>��m��.�[Rcd��$�	�f�'t<�2�c~c؁a;�<����̧�$�Us\l,BKp��;Òɚ����!���|�٥ �~�)U�L�h�(hȮ�O*]�.7?窪9c�bG��@L�	'ږd�5��ω}^)+����l�=�h����3�1�g"����qO��u3�e@D^4�J����?�E�0�`��z}a{�x�,u]��s��>�fC֥F�n� &�c����L�r��Us����i�ZޮT�p�pu`ɯ�����B^��H�ϓ3y��f��?Ǫx��9��u0_�t��Zk��Qg�+c�����B�UƟ�@Yo�0�:�T4W����nZ���������Ň�G^Q���M��N���w<�����|�"�Ed��nӨ�3�����7�F���	a��J��2W��n��Ql��IVl�^�sd�h���s�[��6 ڢ�><.��W�JX��2BX�o�|w���
���GS��������;|\�HF��<�,W󯗣��4���Y.[�{��rM��^��p�%�G(��D@��
xgƜ���_�Z)�
��`���?�	�tv��t���%CD�2��Yh6�U�t��wWQË`t���V��R�y�e���%��x��is?�H!��%�	�Z/���Ga�񍚅��ݓ���X� 4qz�1�F3�7�p{C00��K)�#^�9<���-�(�u�žkD
fڛ�"������
u�.�,���;B�WF�4B*��6��>���j�q����a>jN�$��Y�$�>ske�˺�ڽ5�h{����en���:�������%���J��[�<�o��/���p�\�C
�.����x4숦@F(�z}P_��6�E��UBB����g�J+���0of`�]#iGٖ�÷�1�*^�AV�nBi_I�^�4t�2ل2�!��:>Rs��k�M��b{?�NpW�N_�6]KNF]`���j�EaT%s�V��������v*e2ow�N;�(�<�D�Ȧ����6�K.���ȞėQz�*E�WN��,"Z�.t�r�&{O����W����/�;��%E�^�	�c���k�z�Dn�m"����'E��O���IIlIo�K� ��#�-t&��	��R�2a�`��錰5�䎰0*��Y�tyՋs-stK� c�� �� +j�MZ�}��n��&����d��ǒ���q�q.��`[��PU?h�5�ץ��w�OO�A@BB8����"��I�fg��Ju��Z$t��H�ȅ�Of����#mꈀ�+Qf=��"��b�ǻ:ql���9����;��W��`�ab����P��8�����a�k�Ztn>U:w�����t�f�
�#�#�%7�q�z��c>�����|G�����AxL�����#��w���4��X�e�7�7Wʘ��J9N4?��g�ez���0]!V�* f��.ܿȸ�P���1��Fg(�b�������������¸�7��,�/$j�k@�"B�iJ΃w�Y��ϣg�M�Y�H5�v/�sr󔏽PG�
�|%�����555�d����S�.�y;��Ⱦ�pMbz������y�Tr�T6d�#�vD�n1d���x�����~��K=��u@��G@����OW:'��W��8���鶼���2^0��^��E*:�O�������5��N�;��:R_�n�w��ekzz� G�ᓝ=�t�`��H¡�X��v���@�$J���Wъ��3�I ���?��G����3�G ��ѽ���k�Y�^��U���ɧ[���d%��.N����+�E��ܵ����z=Cs���Y1���d
����Ԇ?3�{K��{�+E�C-Y8�Ϧ=%1H��4���='��xVj�+�u�Z�Y��?,�E'WPh��D�h ,/���"�o���p8��xA^,�� *4�����~2����S����7��T0)F�T,�մ6��큪B`��L�v4 ]Jȹx��Kaw����-��'/����"&���f"�-��g"�k�vII�SC��B�������Ī���a��(��s'#.��0w�n �D� ���.���S�r'
�Lxz����9���U�E3*�E��z��n�Ql^��ej�X{��35�@ ��@������E�.&>������%?��d�l��	˔t�(�7�&�a�c�,��7B��.O� ����NڏM	�N�/LV{"�� X���c>޻�1���5?5�_uR�M����U���dĊ�D����`�w�[u��=`��1��Z>��y������7�5��v�L�$�!2;{�yfNi����XECb���ȑ��.�1%nE��`�R���ꮝi�l�(�\`!��o�&�J�=��5�����6_�ҩn~I�%���ҡ�ǏKy�>
�saoϴ�'�Ya��7���ʉ�B�Y(&my�u�#�M��̝c�d/E������ ����ǥ�x�q$��Z����d������&�����%�[�s�1C��(4�Ŗ�����l|Ve�(�1iLd��3R��8_wtk�AK.�ɴ��8Oѧ���Fj_�u
+�b�3�z�rM�v��������m>��:� 5Y|��F�y�K����hF�鷇�x T��ybT��F�p���=Ӯ�D�S$�ʗb�p?���;8�ʹʹ�Y�O]��.Q���	�Y+��:*�p��< ��R������a�T�Լ��C"�#.��Xt��_��:��\�怦ܤXZ=������lt���5&�L�����c0�&�j���GH�J��;�X@��y` ����^�Ff��Wq  �Ր$��&j	 0���A�[�>+��o��"�OZ��"E{!	��^¹Lo`Tpdxk.ʹ���J��/�@@�2�Xjc�ܚ�P+}�h��[�C��6ٷ2�P�3�N����?;��V���3�[4Q����`H�ٛ�3�hJh�#����?��8�aQ���u ��'M�q���.9���D F��񩩛�R^�њay.������mYi�Dђy]�g:,0ጸl��噘�F1���G�*3*�-���,a	�<T����U7wctѣyW�Ƀ��Q�Y�w���Ĝ�娳-��j��6J��/�*���ռ
1�h"=%,QR8�۰d��i٪�p"#rFRtpjI$(�_I���E�q�Y�e��{���*k�#�$P�Gn�����1�V�k�@��M�9�0�u/�b�� M��
������e��q̕� �Q��<()2����[y�ۈZ�A���b�