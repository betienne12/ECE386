XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$2�`v�`��i�����'��˞���� tbQ�Q��g�]��=%,��&�5��ad�@O�m��'rG�LqI�a�ɯ��up��q��$�T��)@�q)$'��7-|x�l!�dfJ%���� &e{!������������0
h����,7Қ�u�O��g-�&ξ����6!b�:�� {���3��d��M���N$^F��DD�)6����'�:��j57��/Bc��:�]�)�5q�@F�7��xOB�ۨ� B�ԃu��x����G�7t���Q^��3��N��F�Bj�Ca�1Rq��Rd�5�8�pHX� {�nM�7�|G�N��ʐ6/}tZ[��υp?��	��&:�R�������B��h� �*(�NC���F�ܡB�-����wx�y�Y�9j#�Vn5}�O�h|��5a�i֛��MM$�":F����N.��i P�R?(ߧ�0�S�?�o �3!Tvf3���r�i�}k�Gq6qa�TO^�R?�����馷�%�,����󰃸��ׁ"�۔�Z��2�N��#�:l�j�ק�Z��K&�����/K	xL�]'N�����jؼ��~�Ui����*˟���}rصF ��$��<�1؇�0�0�����M�m�)�cgDۯo�H�PB�ü��%l���&�ɾqx���Z��zx�	8��$
r�/�u3��j��}��{�{���xXY'J�����TO�l��SpC���!�WXlxVHYEB    4089     e40����ث��%Z����S���a���װ�^�K��	K{o�S��U�d�d��|O����a�c���KS�? j��o��u��Y��G־p���N�ma>��A�7i�0n�r]9�p&�+���p/H[Զ�_�NϞ��Ct���t��!���y�~N�ܖ�.�h�hc�b��1_{Q*x���؂,�b6����t�$qA;��\,\U�6w&�@�Z[>4 �x�~���f�M�C�=�~����������p�9�K���隌4J�{��a�h�E�Z�ƫ8,y��e��Y�ݎ����A�E�0�`���`�ٴ�n`R�C���{����}}��A(�)�ץY�P�a�OoG*�L؝�q������'ŀ��$UM #U@R�(��j�q �>(QjB�.���EjQ�SLY�`��vc�Bo��]Z[���S�Ƕh]��#zH���Ӂ��G#����lzN�zA�����3'r�=���Di~�e~[E#O��]a��|��U/Z�a��XO�Jj�+RED�֑'��Z��ߠ�z�����X��{��JS,3�K��^��)�ns�C㵐��-��K,�<�O���02\p*%��J9�E���^diL]�?�M+��e��?��g�A��$��r����>D�]<[uE�(���	�.az�1N�+|)+��a�gl���d��,��N��ߴ�ԇ�I�Z[�;jx����R�+o6�@Gɉ�5�ߌ�+r�����]K=S�$H��|YF�#�s��\JM�|���n^ǅqO|'�%�7Ɲ��}(�vÃ[v�,Rgv�&D�ɚ�V�L���3��Z�^������y��1�5���.g��!e���ިW�R���Ŝ��v��f�tw�S�V��{�޵1�cY"d�{>���(�1��ؒ�\���9-�p�i���k���|��ݙH���#���� y)c�uW"��r��r;���w���7�-e�Y=��4�O�[�s�'���M�4Q��i|�ښ1|����}��usd[��V�� �M����ڭ�E���CW�τzawڦ���"��/ha��Ѫ�}�78t�%�V��v�#���S[]���4�,&��1����L_�<�lO�Z¸�:�G@vz&���~��6� R^�H��u�At	%���Z���p��0���8&j8Y+����ǜQw�x��4�v���\�U�)�������+u�?�~	k��.l/�~=�E���9f��w3EWR��M��c�#{�N�
�$��Ḁ,�gi
��
�/�3���?X�KX_&,�a��q�
8�'��h_��ޭu6	[:���:߅���g�-�C�% �.Z�1����99�P��ڮ�2�(�k��ۦE�s���
�d��HMX^���ʴq�x��!��?��']�Xi+i���@Dw�F
��;�f�wRS���p�� 7~��F�M�:4(UC���ji_�1��r���}T<u
����yp���U񤊰���nP)>A�/%9���$�
��
�ǘ߈u�S�;'H��D]W�o)�Fi�s˷YJ6�k�n���3|F0�3��+sY��ᤥ9�pޙ&{��i�ؽ�1��ed�{���ه<����?"j��g�K�!�T'?;9f�o�-�}CHHFps��-(7���ٵ�-����(b3O�mc܄�S}\s�VG?U�&W�jՊ�Ә!B|zSd�L�������ǅ��ڸ�9K�Ii�W�U��ȅ��rz=G}rVʶ���i���Y?c��Q��*�1��eZ���l�O�M�u������a�j$Ȑ��$���j��
E&�����X̒3�ܿ*P�	��isdP�e"O�=J�{9��rz��B���{oo�������(0��d����_  ��
>,�r�VQ�x�#���v~\���u��\X�|ݘ�+6'Ԙ���,�}�4%B��3[�.��S���v�r"7n�6p8��L��@��	&�$2o?$�o��t+rjɥy�8�N⿡!gh�#�)�"1��w�œR�lX�0�!�:��G<����"m4�&�����}�t�#�hk2�]�ȜP�@*F�\y:�l�R5y�%�L��iΚ1�Z�5׍���$x��MM��ہ��ڌ�W8s֗��2�L��+U!p��g'X~֛�Xm(چ;`�׮E�@�!���!W�7RF�V��U���<�ӑO��`��Tj���ok�^UX����{����T�!t�D�T�[�t�������}G���/ػ�&%��i��J8+�f�;*���0�^�%8��\��1
wN�kO������R���%ha�R�\ˋR�8:��㦰<�!O
�0�Vz[�pj&��	�����WD�l�k�$���tG��Ǖ���~��/1Y�0N�a��h�T��YO�
pbNJ~��Hl�3��S- ׈�i��p�nP�9��m��c��7�N���/���!��S�0�ء7R����"��I�^|vN�+��=��$T7�ǵw'�G1��"������<��`���xc5�:YL9���Z��Oԕp�������;�����lE�R:籺�_��O��w���۰�[�D�����3��1���l.lȊ������]��_���J��?�w�8߳����i6e�Z
[g���rP��|1�
R9?��m��������i�~Y-�<���
���q��A^�U�>$*ͦ�g"+l-�����+O"�;����[5�rahX�=�Vq�������Foa4
T�-f����5��,1&�������������o�E�Q;5��B�E��K;'́�R�F5�kd)�\�K!mNc��+%Y��f;�h#f��#�S����/�5y�2�s �"��ݩ2�-����y;�q02b��h�8�]َM]Ek%ov�oqfc�\X�vG����cT�n_��g���n�&e�Os�[���ַ�Ȳ��1��1�(�B�p��a�f�w�aUҶ	֬W��g%N��3���n_�2R�^|�r��XԆ��8f�?�����$ �k��6d|���x���b=W��(|����~Un��qI��d:80;d��9�K0oQ�{�&ˮ���_��ˀ��8�v���M�duZv᠆��}�6�%1��́�F�2�X5���ڶ7�uA
��Ɯ�W���p�+=�H��إ��21�^�ΒCap�B��$��h��`&�b�vn����>f�cI��0�b��8`�`��U�ݬ��A�.s�x��A ��z>�x	��=qy6R�Tk�ը�A /�և`�e�y�̯����);Ha�>�?��e-!��+���W��s��.<mz�0��BB�'��a�RD�"���ɠ3D����J}�̚���ݓO�|�3��t�݌��!(H%���j���=�Z�l�:������1v�K�<}J��`�����9��"P� B��v���e-�i��Nj��yW�g#���1�Լ�`�8#Վ&�* X[֤�z�S՜;��g�G)�6�n����ǡ6�? N����^��u"�\�5�YqR�������cl����a�|<�`��7^��&�ƹv�ÿ�Ϳ�n�ғl�}Z�R!�a,�m�W��SϓA(s8"