XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/�fr��k=GN�6�y$T��g �	i�r%W6����Ï���/�!E�q�m�i���E��6ƏmD��\��9N�@������!�voSi�����J�SC�#�7<���msA̴�y0l�.�wB��2�u:G��� �v�I4������/@]U�sR�0�<�7�' ���wH\�L	��}tau�(�~���7��i�8Q����*C)i��S�#����єMã�2�t�k�	�r�"#�j��z��!��^��Cb�EJ�@�5��]m��-.V9��m��P[�7�s�S�Z�mU4&E|��0��¢B��8
`����ș֜Y�ֹךl慿H"�SW^�ZTj`�U(��g���-[��5.�Wr�P;p-&,(�y�'����t�&�..�a�1*��4�wϠ�S�&[י�E�*�C�j���-�s�Ġ���JQ��Ab7�F��N��\ޔ�!�5~ʯ�I����K^~�e�%� �
�Z�	�)�6�ٯ�1�'���Iz<�'���'�P@,U�&w���Ӆ���^��[Z�+p�H���I������-R��G����m�)92����+�i����8|| m�j����V�gf
7��I�	o.��'�$H�n(��Lml�����&A��s���*����b����2o!�8$�%3�6b���/8�&^���cn���zC2H�|[���������^�,�������dǤ��P�uZya���f(�Z�~XlxVHYEB    fa00    2470��:�jP:�1'�A�"
�4'�W}6!*mV6�X�N �P�
�6�_�]q�<w�K�~�BI�.����>�3������/�k���N�%�J�;$n'L|�Z��z!c)>܂ ��`:�����&��H�|@��S(p�ZaԱ�c]�fP�I��L]l�,ǃ!�s�"��\o��送��XHC���Ϸ;�%f;���~�P0�g>6G ��u'e9w��`%�;�ӛ�^�gm-�N�$p[ջ��C{.CS1�de� ���L���8B��|���pk���a!R����9��-�Վ����K}@��iAb5�������̙�ΗB�ec�5|w�sO�+'�݌�tsB�ɺo�:�eH�`DG�{`�!Т�q9#A�9x�~�8���$���E2:��sE������9���w�]�г�ڣ�Z�hw��u��B]��sB����|\
��/k�X���2��>�ה�����iN��y���b;Ē�2#7�c�Q,&Y	X����b.����Bdu����t��ۚ%�L=H�����3�T���t3XE��-7�+��pVr�p���@���0��v\�Z9�+z"_Q?}�5`�D��Iŏl�=��*��xo�����:� t!W~�V-r;b�ZJ௔:rK�,�4HJG��#��J�����K�ma��b",��v8��[��J�έ9��4��#��kb�$
�E��=�����+�x���_${ �����I�_&��)���w����e�f6<�~����t�"�g���P�<�2�����g����H��L�}��+ڗ�K�U)��~�� ����^Ӗ|��9��S�M�]�`��0���U��i�u7��Kw��@�E�C�%��֤R�ȿ���I) �����N؄f�68���Ϭ��6���K��BC�գ�a����E����H�>V�F^a��2g���1�q�*����f��k��/Z��v�;����^���W��L�+�>,�3�:�^��Kls�r�(�-���φ�bc�����݀��������c�|��	o�Z�xAuf�
��&���r�+���b��Eմ�.���<��ѻ�����`�i�����$�S*ΘtrR�|Uc���pZ܈�����L8�GM�l����^�FT��8倫2�%�%�h�ʊ5��2�>V���l�$m�e�>$�~G{��Ӷ��_\���W �b��#�P�)���-����+p����10_�"�i�;w�.l��L?�2r�&��Q'�y��..�-���hO��b�/���!�u]-������7�!�7{.r
�
Di.�1��CHBҢPbW.��|�/�i�69d���� e�As�Y[F6�i��-.*�����T��_�}��0����o\�J�dv���Lj^�H�d!9p7e���v�[rh�M��{t���*�����sAE��+Q���P�t�c\5�,mꓚ�B1��z�������}��#ժ���e:3�Qn�Ϩu��C�������������1ћ�����O*�Yq]ަ[ �ƭ�g����J9�Z��,��~ ,���n����{ ��ϻw��v��5��#��bqRQ��]c�%�<
n�>sa#���k-�W6Y_Jl�?vű�@�~�/�'�O�
���R��Jk:�c�t�i.g����\�VC�����}�9�M-��VJ��T�����>���ܵ�'�^a��:G��z���b�8���V�~����'|({1z��;�dE�
<��2��L�\�0������p��~2*jВ�tަ˰뗜XRE�3����� �8;T,|�'�9�����}��L�F�ꌛ����=ΜDS���dԵ<B�/�D�Oi���J�{H�9I-L�[��/��x����A�F�,���%��#@6w��\q?��T�H��E��O���g���mG�^@K��^"����e3?�����s��Kl(�TM���)M�a�d?�'v6.y�|��^��0�z��i�58(Ɇ���x9���u�]�-6.�1S}>��!d���g�l^�l�t/=��/�`G٧����$������~;���Z�[�Hwp�S q�[hb�@c�-"�p�4�i�g���1`��YS{z/6K���N/e/�XvQ�;;\]����X�[Ȃw�4A�Il)�������%`Ҍ'�l����@[`��z�ȟڟ �d鷵�u��7�.oF�xFaŴ�v��Vo���{���WiR���kX�l�j�z���F�{9Tgs]�Վ�����d ��@2�� ��)A�V�96�rT�i�6���R�-��8L�V8W��5qv�u%V��^���
e����2���奵/���)G���x�&{BL�$��E~Va2Ѻ���ES�dH4�sU��wE�J�h�*����JD���������sQb��;9�����s{r>vH��E�$!�-@�"h�p:�-�W���������1'�jZ�w�~��)['� ΝJ�cc��2@�V�� ��_ݪh9$�|��Kz�"|�qW��}-�vĆM�T�L����攐���
,v�*��D�5X)X�s=���Bn=��44�1�+����QZA�aL���
���>Kʙ�����u0B�+����*l��L�����8gM�z JY��A;"�A-?������uDwD�'��	g&� ®;"�.��P�Nd�YJ��
�I�$_� �T�'�~�D9��@0��L�&\��^��%8̑U�g���T����o���]Y�e@*&�zcw}����&�����3L������<�YҘ֐��<"���;�6���̕�K��ϛ��9�ͻ��r׵���j���kX^9���R�:1sbǇb�,��E���~G&a�m�E`g<��j��7Y��jF�E�H�R�p��f�6i����#�0��H6��<l(B�㊴r��Pg������\�Ӄ�{������'���]cq�5$9�^G6�x���d�o��POِDH����k����D^UP��ݢ
%����(�=�Rn����`�-�D����u� �RǙ�b��ܚ��s�4��Q�<�5����w����������0��8�d��\I�A5��gL��sF�L���Qtڝ��x�6f�P=���rwA�5�	�Րz�t?*��K �n&�
:������s
��"M1�C���)��ݗ����� ���9��ֻ�5e?��}��/V��c��*RlEa�ւ��B�dj���~��$�G���P*gY�l�d<~�;7��ۀ���H�s��2H8%n_�V{F�*I��0h�-�1�w&UN�k	u���s�U�vk��YP���[tD�c�"0�U�Z��ЇB�wl(�9��x ���p���Z)	i�Q7��@��P�.~��(~׃�ͤ�Sd(�>��h�h(i ?{����Y��m�<�'a�����E%	at�u��+�9zn��<�N_N=&�� �.J �f|ʚ���l���}j�6 �����,º[DǳSf3g�"*|�'F��N��.��t�q��E\��X'B��y�m��z�\�=|ݤ�<���;�?Q _��$� ٶ���aǀa^�I/|V����ȉ���-�f贉^�ZXv��I����7�C4�L����w2���OǛT�N9A+���26����F.z�09�1��5[��F�F���k�m�/�b� ���u=�	�#6��v�z��sd��\*�Ãu
׻�i���u	���r���&<~�����I_P/��9�\����k�D�֞;;�~�T�H���/L�gasY�;|�[+����'���������:�Q��B�IX��F<�"��8����jN��rx7s|J�����
0L�`1�6�͢�\Xm����������1`����J��e}����<�ث�ƆQ��>�p�\�m63�Cȼ奾�B�p>�45i�%6�FXCr�u5�&??�͏���pw����j ��	�w�1":����rX����@ě��4�|ZuÂ+��S�v���l.������+�	V{��k��{[wz�nyŦ�PB�)����?�Y�3Rʪ>����6�I�o7,�����$��-)�'���bt�׷+�-�ƫ���wm�晥� }�Ԛ�t���㦡�&�IW�zs5�X9W�K\0��6����°��
Cx��_kMöL������P�ȴ!� �������j�01�H�Q��h��>�)w�d�`q��]��,SUU������k:o5`�yʾ����^�Q��\u�܈��$�m��[�I���(2p���E�%����z��jC����L�^���b-��`w�F7�6�dk�p���l)�)��Ai�5������
 ��{��Sa�����` �)]�WEȱ?Nq��3��K�<��ǽ�L�^Y�[� t\�&�6w���F��J{�,��m�[��,Y���<I��J�f�S4V5��Js�s���n�Ŗ��)�OǨ��2�G���wu�t�/^�3A��Vl�ƚEѤ�ͽ���j��՛=%���9T5�`�e��f���{h�B���~���$��O:��_�+JP�_f�u���Kg����[՘<r���&�H�����˜X��
臓"D��_"~�7>t�/x��ĳ��L��>v!�hoJa0��b�aQ]���y�,�u�Z�ꖐ=�*a ex��Ul+����Ɖ�M���`᎜��e�w^=%C��"�F�·A���pӛ�3I�[Y�A�Vx@�t�/T�B����N��[Dk �i�\�.h��ӛ�Xp������K�����!nx~��b�g��,��������)��u�A����ږ CYo�ױ:��9�F�1��~�^q��7��^b���UA���C�bB�6��(�+���(e�q���*7I�a�b��Fg�M�7�@�Ϝ}A��>�]�9���#��*�<�͵i͈FZqbɟ��ܐ'%'/���7�6��ĉ�pz��)�@���k9}1��&7���f��*Qb�h��F�~`�.� 	�;�N�
K�M�	J��;	���>�i7o
؟������޲*u �"-M��5�&�R���1��)�4=�e�����n����L����N��)�xy譧ܪ�1�3�ܛ!Ub��Z��Vb�ӑjB�}`��n<�-νXC2 ��h)��ڼ��#�|��o7�t?t<(0�������vaA��f=C�zK_��`��a~Hxe!�W(9Ө��	L�z8�;�_kBh���H1��1)r��%���ɠ�dȢ��u4S�0����Qr�	5��bKƘ�4#�P��%���%�h$��� ��z��>�"f�P�=��_���h�N�����x�{y�C�jT�FE�Iv!m��������@x��B�h���S�2 v��)-��2�I��vG����Ni�9�����ّQ��8�d?KX7ث��ۍ��"���>9�(�&��5x����vf���twB����Nq�0�-wE�7!i���3ۇ5�L���$�
� z>X1����Pf���͗��m]�g$ ���T���������7��q���E«�n�~�f��`�E�7zt�e��@Q��豮�$wh�$:����|�$)%ܙ�ḋW_lN����q������փ�IQ>��
6����bn��>�K��(�[���}���*֯�P%��qm�Қ���&*D�̂���C���?��_Ǉs	��H�Y�K��O��j�C�,�@��ދe��e@��ӲDz�m�$�����%<��N6%&�Y��Pa���v�%���Bn�go���Cc�T�	b�d���47r���r_��gr6>""����?`X�ڔe��Y8�^�����ݰ?�U��d-��c��N�Z�"�;�	p �z���d���{�+yE�]��&�Ʒ>r@�0m�k�م7Kj����=��x̖{J�p��mA�̨��y�!�?���z؂��4�u�y��Ts�iJm+X�D��ۦC�ئf)*EU/,(v�5h�V����#T��\��|��S���L_s�>1�����@�7�K�?�g�U ��{��|7��־�:�ϝ���N�&Jh�\m4���.�JQl4�VfN���*�r��E�ً|�5�ѯ�K���7%��mg IZ6 �C��S&���
I��Ɛ�MDA��?!�2T�V8�c�0�q��b�B��%�J��n����'{6�pf5%B$�^�=&G���8;�*_���F !X^/�)ᕑ��1=Uw-Sp)P��L�)���LI��-G5�		5U)O��At"0|�
�;m��y����-�k&�l��
�И_�IK�+q�-�G�ob�k��O]M�Qs�2~�ɤ����SN)͹������%�~�<�	�!eU@ �귝G���#��#�Sw��[3>�՗99�ߖ��ܿm#��@U7X����{0n��E:f2��@���zf��	�Dqh�_m-�]�sի�>E^P+?��S�t�#��ښ������Aw���h. ������@ڠ���꼓�H��a�����kUS���XA�8{oC�
���%lgYy�����wZ�nP]��K�D���u�vh�=��n����_�b'��/5ݢM�n�7t���,�Ef�Ю��x�l#��G�aD��#�5o�V\B<�jf�-�w���d�ʥ#�=5��9�FĞ<�7~��H����j6�?�bNBA#f.oi����uy�g�2�{�$�V�,���!7㻣KB_ǘ:�3\�	zh;o�W��#/�li�:"�P�s�!4�tt=y"�UR�����޲u�g9�p�����-->��o���m��n�Ů#�R��IFEڼ�?����|��SO��/	O�����e��~Dn�O�U�
Q�&�xy����(��	�x�қ�}*�9aBD=���u�!���p� �=��TXDKI�D-��'�|_���x�5}����k���%�ȋ���@Q�`�t��ct]c�J���D�J,��K�(���X}VC�å=a8�AcC�\��?o3��C�h����t!_��=�t�ӛū>��C��*�h�Slʤ�1��7v����Ls����J�CU�+���>/W+��g�a���U⩼uhm}{Y���8�2���-����D��o�Ӌ&�IܓG�z�T�	�B��eT�X�߰}�M'pq`Z(ZpZ�5,��{[��0\�(�v�r��Dp?x&�B�4G؆*���t�S�*~�P�2�&�cb%
���VzH=JI�F;��8�� .rɵ>����~��d��Wz�h�2k�=� x����Mv�xH����U߁+��rP�S'�~u��@��Ny4������(�Wj��i���,_�*����1F2�|��lf��ۭ�S�;ŷ&��C��ƁdJ�O|6��Qˁ�AL�4i��!����D�Es>��ԇ@���`
��֛h6PE���}F*xT"��R@�c��-�Z�ӟ['�\�m����J�[/�W0�}�ʬ&�����(�u(��j��5
m��P\��X�ȟ��U�=� �K�;�9/X��3�]J ,���*�$���d�yYZ(�O��횱L�21�g9�nP@��Gy����I���d.F�V&��H�zb��ML�x��+����Hkn�iF:�o(P�^t���������$��<�˵�3R2Us�o��2�M�Rz>��j���!��,=5���/�=��4?<
�q�� g5�-~��_�y����t�N�����V�~7�.\)���k���'&������w՘ʻ�������԰r6��R)S2(�q�.v��{MO�D�Y��>��p4 T���	�Ym���?�
��AIC���JxSfN�A�����}X�H ��H�2�z�+]y�����-��&Z����\�|QQe-���rbp�)�웥���.:�U:D�;�s==��.��aB���Ib[]����es���K�i�К2�]a�Z��n���,l� �K}3��Tm�u]5(�1�{	3���|lwP������O�� ��2b�4�_��}g��!��9W^����ͮG�5%�#Z�JK���Ҥ��uC��$,.��ir�ۮ�U:�����A�B���?R��F��-.��Db�p���{Z|��&�~�|�~ZMܿ���8����d��䧠[�J��a�@ȓ'6lC[�Kc��6:��ǘ2��&�����ZWϰƿ�G���^����r�"�q�Wn� ڨ��i��f�u��f~�e�RP5M#�ND�-�)h,yz�_"i�?*yf�t}5�>�)vʏ�?��|I(#z-|���pa_,�֘h�f=���d'7�r���J8C��ʚ�e.���.�i�ӿ韘��2h4Y0I`
l'�N*7B/���B�C�Z�G�� d	�{�y0#D%��Qyw����Zj�����%�/�w� ��fS��*�]���~���;֔�t�҈ ��h��/�}O����|G���>h@�tȕ�I�5MF��a�LcN� �Y��2����[��%^J2�|B��w�`�����)��(%�Ф�Pf�K*J�����<�˧�6SA�K�yU��~���3��뉀M#�Ǚ(���&٧k��3e7^/�Q ���מ�r�o��u�!ru\�U(�~fix����ĵN�l<��+&�^N�W��o��.�^V�5�x���_u{ª/1|����>�+��f�4F'����[C�
��M)y����ޙN�!��3��}�d�uݳ�έq"qB:��b�f"����e��'t�����Fβ��,&�.~��Bj�p/*��zrڨXF�Ν/��4|?L�2�{�M��A�PG\�m1�>�B�7����YOQ3��p�)-D)��hN�-�QI�&��/�W���<Rì�3�vr:R#��}}�=���I5V/�.D	�'���͜��NvR:|��e����h9�&��x8C~62��9(w����������"�?�c������6���9�Q��+�����
�����K[��h���	�bY0�����$ŴI�Xr*X2F�걬����^k���$��q~�IﴑLDK�M��UƳ&l�(��)�x�A=݄xb�"���[�Br���~��U��[��,0��ײ~���-�HXlxVHYEB    fa00    1b30�6����M�g�y����7fRZ����e�3���i����#���2*�q��}K�}��Z�����_��"�|��]�^����vm��5�X6 b�A]�t�<�,h�Ѝ�DQ�A?K�(L43y�:0A�f H}roB�B�"o��r풉^r�mx���H-��/��\l�t����`��1�7�\��ԴD�A{��6�w��Q��0�Vv+.�h�}H�mh
�'K�����HU����n��5Sf_�R�毞��ծQ%�= �������m	��7�%?�y'�S�:U��w��9�ZaNǈ����W+�w���<Z�J���|]��f~`s����GED)��%C��n���P��^�������=v��Ѿf0ܡ5G�OG��oe�Sw�C�g���XDz z0펭?Q�.th晆��ZB7�i"�j�|l��+�H���ᜣگ�7,�{��Ʈ��VF�q�<�3����]�ݡ����f��ߪvߞz�����0�Ρ��/����-!���̣
�h+lQ-��!_�{��hR����`X"Ψ/ͯw@�S(��$Okt�>3�֟�����|Q4Rb1�TB�ᮀ��Ȇ����5فm�͘�u�����~�o���F���c$��#q�@%к7���'1��m����P �y^�QOw�!f	���^<!Ī������
���A�����h�f���X"q	���dDn����5����w`�a�9�~�o��
�_5��D���3���v]?���N���|�ί�k����5'J�`���}J���[��b�|"�p��݀�J伔	�[������	�qFh���G/o�t>p/�c�װ�r�٘}M3ΓNep�w	�������)�{�Z9���u�_�T�ފ������ٴ	ۓ��f�V-g=vS�}b���^3�7+���_�����B�c�\��8�&�%�A��)Ey�%4;��z,A�o�+�@V*��A�d�=k���:��]����yǯH5�ҙ7^n���ظAuҭ�$+�?�r#k�8�����g��e���@����8�b /��`09����B�* �$��%f(g����"c�*��Gb(����?�)��9�g�Uvm��y�l"볱i��r�=դ�~"(�9��h�߲�¨��M�̗Y���0Tf���$���:���2zZY X`۪&(C���J�k��#�F�#�-)ssF3��j��?-ą �(Gɒ=K9��{��n��l`��2t祫U����x��[���k�gz�=��r19�K;9ǈ�z����O��6
��v��� �u�:֡ob��P����D��YֵY��W�FXʶ6����~@�N.��ǸԌ^~�Ҽ���r�)����$ߨ���+[WK;:���0	�";�Q�5ř?f���;p8Kw����E�I��zv_BL� ��5&��_��#�<C%��>�p�����)�ǡ�t����C(�O��*�5��NB��CO�!`��忁���m�\M,�WEφ���/>���%�5X	�R����a��a��(�.u�Uz,���ٛq-)�K˒��on�u���A7��s	���;3�����n�;��jC-�x9Ţ'�Q�њOxb�>����=c��Sf���._K�u�B5��!'{�%T�!�����_�RZc�!�����TLg�k;R&KNu����@�q�2�E��
f����l&�27_쉆���5kQ��/m�q��$!A%	��8u�����j���j/�`�3-�T�R�0�AVֱ�ͪ�h�w���_��ϜZ���9�۹��n ��uD�(�!l�1���F��J��'�r��� N�>�V��1�����/�-�l��8P��д0eIsS8W��>#�����E����v��߫�:��)z����i��d�_U��R��.c���Hv��Ɯ����;�*��8�+Q&���t�,�8�[���6q����e��kh�W�B:{~]@W��k������������@4�ߤ�}.�M���db��%	��S�� �w큯��W���·�KG}"d~��[%jn�w��5 �m�h	%\j��~�w�8��Ҍ����)h�bn�Լ�=1f*������Rjs̈[�#��&����.O��[�pu�K�e8�ۺmy�3>���KJ�h��n��\]�
���.P��
S��������Qm�� ��� :��yK�8&i7�?и��z#��<��(r�
�1��Bp$��D���D?1@�(ݎ��%�O����m�$��T��Po�iq��׉+�d�zm�F�TPTP���U��z�ί��$퍵W-���u�rp��tըy�_�Gp�t��r- ��v�}:(����%��  �o�!hEr��>o�,���R�GMF�O�!m������Q|_�j*Ჾ�@�ю��x��4�甦��>D��U���8��2������:Q�]oE�r�i[8������\4T>7d�r���Y!dl����`4�v�@�U��8���H��n�S�׆���W����~��MI��=<�L1yگ2X[0k�1p�֚�Nu����<�uJ�?�z��!�wx�����U��C��mz�m���rNf&�AI� ,r�j���+������Vcɣ2D�n�̭��P�#��4��?�������N�.�R/�?+�
�ጿf��m��i�Sd��2�eQ�8�Ѱ�G�{�x��wB(����Z)q/Q@����򇾹O�=<)E��u/+� i��h�)�=��TU�p�. �"
�+�hK�WC�nA��]PSW�w��%���5�*�T-:&������kv%��!��[�]�[��jGaY�n����A�8�����=�8�'�n�JB�_w�3�l�4fe�i(gB��缟"H�ޔ��f<���LJ{�݊�͘�ښb�Ȩ�5e��c7L��x�O)<�Ib���#WZ�Wo��	�D��	��j���0Pj%I����J�a�\ֈT|���O;�f��f�Q\�>��[�H4_�1S��a�|�))�I����Aib�=4r�F{t��UK��}q`��G�8����<����5g��%� y�RD�Io섺��F�g�qk��'Y蒍�@�{���o�q���{
�l�J�K��	�6K�ݤ��~ sɾ>���}��a
�x��N��,��MI�4���]�`cfÂ�b-Ƞ����zBvâ�ԗ@ȉ1Gq?�������O�yP@1Kn(jj��"W�0k��Y�.�\��p�7�r��|L�+,L>_3T}��p��U�r]��oT	p���0��}�[���-��8�xx�A-�iLK�w��"�������z>װ�di���`<A3*��W5�Fy��jMW���2�}T�HKt<�q�W���.x�s���+B��A���������.wY��
��Q}�ā��o;80&�q�oqoW�X�^��T��9.�A%>��-lF�L��-R�f質���9��k�:ä�I=nE:t�c�3�|T�c��k���ݥړ�G-�����T��i�kr�
�Ō�
*�,Ya�������UH:�Z��� ��) ���+��B�B��qs���aABe�<�)y�
e�E6�/sW簧M���o�|s��ٰ�����!���i3 �p�9�P�%[^��m��ʐ׵�~$9�O]� �W���70/"~���0���OU|t���l`#����O�r_4�[fG�
�Α�,�)� 䆋6H��H�E!&��w�����G��㳜�ʛd)t����W��,��	�=p��I�Lsd�2��icXJ�CU�K�+����T��Ad�����p�i�$+���g��[��-Ш��[Գ>���]�$g����3�7�쥰���$���8�Ki��=<{���ځD����Յ.� Z���${�_f2pnKĈF��ha�-ujRc�r��n��f,k{�W�E�3�!����έ\au����Ó�2KaC{xJ�S�u̦�c����t!T� bh ��a�;�z��+��[�(������L���CB*e���8c�c��a����e�#iX6V�pq=L˅\�E$��wɯ����j���|_�R���E�$�o�r��[�p��P#�E^j�)b��_���mq�����=Ŵxq�	rx>T�
N����}%�yB ٕx�J63T��D'�Ƙ�ܔ�"��\�Hh�4y���*��} :��3-��߮	PJ����� e �������b�y�o�7.��[�+�2-"4E�4�_�{xB����f��\h~D/,1�ə��y�6��A��x���3�C���ZZf���y�"��e߿�?)m��A�m�Ul'���̄�ʏF�l%�LMl^�?n���*Ǉ�%[�H��x��J�2�����u�Sr�(�<���mOb�!���G�\3G���fs�� ��Y�?�w�T]�,U	&;�D"��uB������0�S�N�Y}l踨0��}��q$Y�Ъ�.k�` ��Y��~��9)u7�"J@�s������f�x
wr:�{����a0 ���ah�}�SE_�W�����~ ݁�wm}Ձ��+����$!tD��:'m-���u~ Y!�O�C���/���$�Fw��E�&P� �Y���.���L��kyZ���/�������+��9x����|T���Q��"��6s6Y}�{e�:rTx~^�IҗJ�.>]�.%;`٣���2���vǁ���[0X$�(ْ����T��~�6�ʋ}�@��=G�G�Q��s�v�ۦ6�l1��ה�EJ<h�{2O������2��6�#���"E�	�K�$E��`B_p��Jw��`��*�կo;oɼ��8y(xu�5vP�m=�*S���y��u冠�7�8A�N�����GO�K��O�����9���?�M{Qu!�E�I|T\x�0��j.4L�FAj[��p�ׄB�\&b���/�BfF6�M`}�|�a(_{D+i�������m��`����x�Ff�^�(D_�:�@A���O�F���|u6�lt��uv����TKitնO��!�a��P��J��iN�q<k.�*b%;�&�̎��2������y���h�kU�HL��� }=���"$��	Q�j�ngJ7h~���~��׸�8$���1Op�b�!k
}	�% ����8u��7+���,
��Z����0B�;��So� ���<i�����F�ܝʷ�t[ߏ�&e�����y�G�kO��9�Ж���.iz���^=�2s�~��Ɓ�먤Ǧj��
�-�<��>]���졿���؟�b�&eo��ʢ��5˦Dx�4�r��\:��4�sH-��
>|��EuAnŜ�}�w;�,K�NM8&�ߔ���aE���c�or���1)h��i����G`��:ʫ��3]�P���[��K��^ɵ��t��cΨ��=:�K�#��ȱh䀱��t.b��'������F<����� ��^�:��v�D���9�.�<�81m,iх�T8���{���z�|�O��R_E�5��X����J���{�g�����.�=ěbz
�Ƅۮ��,�d���pu����;M$��b��w'������ ��JABr:1*9�����*�a6�=��d�6��]զO��a�s� ,�2hq�:�F��!Q�~E��ml�g����<����`�a�ḥ	�*iPv
�T��oNm�K�G@��w��c#�c�J�Fn֒�[����"6�ћ�{��b롣���O餷�&��f����E��i��RE���#�OYE��7%���z�Zշ�Wf�Ƭ�Qa�P�Nj�X_%琡��֚S����P*�`'%��F��f�|&T���\��pAN�fّ2�M�մ���p�� }l�[T;oڽ!��~T�=Y
�Q�m����;z-�_�c�6;D���Y��E*�R"��D�]��Vu���"0AA��O�����m9,�<��Χ��2�S��:��aO�%��U���\��N��y� |Cg72:=+�.��\������r���cƖ�)X%p�J��``�"�Z��iop?t'�a�B�Ğ.hT8�;�u�7�%Tۄ{@パXt�ɷ����z`��o2H�2.�f_'x~�ƉǤHUe��"u��FS�V�ZA���V���S\��v-s"�K�z��s Uѡd9Z����8�qn���j|������F�o�c<	���	�GF��S�͆ƾ1y{嗜.qk�;�@��s�pf�t�D��֨�7]����~4 �1��gs
֮`�2�˩j7�&�<���%�jѻ���^�������9�pN���sբp2���ԹH��9`a�QI�;i8A�%s}����Df�e	hR�缂1��[�&`������l��Y#�-ѧ5��
��V�6֤ZP�Q2�X��ǐ�}�&xL�\�	ǿ��%�x,lnI��W��f�m<�>+���Q�R!�k��o94.{֨�8߄�� 0�Jiy��7�U���8�E �!+/��IK�#I�]�L(?L6FJ��6UqE*�\{I$�e�gbb��T� �����1���̝��P�ây����Th����+���s�e^���X�`������a���ۏ���noaӽ�\A�s��S�x�[uM�6�,���ѾebiR�4�51���Z0��=�~:c��v��!mA��h}c�:Q��
)�7Yv�u5��c)����l�g��,�0�c\
=e�7=N�<g�u��aykt�j�3�U��rWC������%� L04X��.|��>Ϸa��� R�z��6��[��C��5dH��|�OXlxVHYEB    fa00    1950`�F*��U�I)K�4
6ar�7����ͱ2��8'��y,b*�t1E��t+�\��-�6�>MهP	׃O��������DH�����Sm/��A;�lm�xV�]vY7?�LQK�9w,�	"W��e��v���^��{d��e���)��h��X3�rV�s��SmL-"��	�f1H�M��G(�&B�;��(�P��KsTH�<���4��>+�e`�⯨��u�& ��TE������	�Mz������$�OM�+U��,o��pC��b-�&�ӇDJe ��ǕNed�O$�l�E�Ω=�C��y�(�E����g�O�0�͛�G^��I!&���U����I4�b$�?\�XV�kE5��
�&>Pj��2�'���E�Ο�P�-��{����}^Q?ڴf���~�4=��D��<5`���7�-W�}!�����(�b�!b����ډ�/�y0?��;K���I`�;����U0��(�����
�汩�zv���*��TGd�6�E^��U��WMR������m�:'���ƕ����'��g�B�2�[��&�n/��d	{d�̏��u4p�=�׎���{�K�7�[�B�:��g|0�ݟ��K��>�Y����4������}�	���dRY���+����+�`�!`fE.�i����>�w����[%pO�!�&�Ea~uN-#h<`���Or�p|����C���Y��@'���.@øRHP�(ޮ�jD��Ҿ�)�t�)��.�C���)3���S�Α��/�_�(!��Jj��h�J@��7*Խz� 9ڧl�F�@M-H�'�9k�әS+|k�{䊗�UC{\I'��7l�C�i��fd-]>�%N�9iX�����ӽ�e]T'<����R�O�?�~����0X��K/^�����|+Ure�)�^�D���7����ձK*��&|+Z��Jձ�Z�l���7�!��7�x ���5ڑs�,��+��w�#�/��ӋT���A�~U��E��ZP]��{�gk�;���mR ��xC�����7܊ ���t�a�KR�EcEA�#}m됩����=VK�4 #O��p���3F��`��� Q��j{�A\�$�!���P�
��۬p�9��]���r�I����Ϭ�à|����S��v��>�'�3���M��IGao��@���3�P�RH˲�kN����,��$�:����a3�QK>�_
8J�"�ccK(�u%1���YT@x��Sb�j9yz�*O�Y��aĂ	�$w���J������ŝ&����T9!CJ��j/G�l��M�l��}��8.�M���־�C�ݫ�]h�d{%�P���.���av�V�>ɄÉN�"�8ܞ?��y��X/���)���e���	p,�	8c�!��-#��� l��Cr��V��#��}{����IU�<�霮r{+;�<9�V��t�������0\����}�wWCة�V�3{�d��;�ƿM4�kI�b��#1�!2T� ܰLd����vś�k�-R��)��Ra���t��'fXO�H��������n�a�qd��]���J�>?�D���j�����~_2��Ɨ�ks�̯i�Z.p�=>�b&/c�6u�/<6�|Fؿ��YTh�ߙt�V�L�����߆�9['�:#Q�;Q������lvС����K֟]0�+��|���T����v��qD�yze���G�}����N�k_��@�~��FI���ˁ�7�7�O��©8:���>�X�_m�n<ڳ�6j��j�e�,����Q��v^^DOF� �'���~o��~��Wz�e�QWD���t�� ����N[���u�����Tp�7�^�j���_��=�+S���rr��,��<�VGti9�7��/o��j~w?s�� /�
�~}�!��x��[�qhN�}��?�;���7e��'�:ej��#�oH_r�� [E�7�,k���4�� ��Liy��O��`�RT�s�Ij�Js��n6�_~;��H��VC)�OX���۩�b+��3�ȣ,n��]�b�D˕����(�m?٧�9x�h�v=~"꒨<��2T{�z��s<3�Gj�Gr���5L�3J��$��1�!vl�»:�(�s�.�kǊ/� `����J���}������ݵ�'J�j��T`C��9�v�7i���U���^Ϳ6"�����
��t��LpXfR83V��f<>�5|'�:�{���$���y��j��wZ��Î�� C�*|��訓�)ǫ]��҇7y���iT�����k7���UY�)g$p�i�v*�kAѻ�rD��� Iw��NSǝ�
�w`Z���HQ&���
 :p�.������Ab�f=v�A<8ZI߇M+�vFa�+����X��ת���9*w�g�"i�&��Nv�( TPɔs�VW]q!2z���E$��!$�L��^��{?�Y��2ލp��2i��Q��=�jq:^��~pn�!$3��Ф��c�������#�d0��R�`E6���v��}�TN�MX��OI��ZYs���T�"��	�8�w+k���w\X�4�s��a���񤬷kI�?w��in��[�F�F� ��`եhǰ,k�����~�H��d6^��t�Ĝ$�:�>���e�.���ڟ>�q�-�?b�A!����Gi%&�`%<�ޙDu���fd����R��\���Cl.a��j��r�g����.������H��Y�a7_K@�ޜ{$@�޼?&��¼�E��l�u�xW���XZӦ~(K�;p�[i����tf�*��g�N�������UJ]���Uq0��u��'��vf�.yWM���L �.a�+�P��L����/w�@L���3%F,ٸ��̀��TZf*��R8�{�i��5[���2���#�2`��\�Q]y�Ė0�Z(L�L�
�^L�(lE>��1p��7��3w�S��E+������ǫ�2�n��iMu���#W��*��S0C\��T<�.ۋ�kgy�\�vM�ϊ2@��n2�j��x0rCh�]���s�f��)������L���~��6�7"UA���fANB�e�JO�Q@d��,����X9��W<�h�z���;#�u��ႁ��@u�c@c~-���m>H��vkM����7!$!C�IJ� ��g�ߪ;��~��kh�st8nߞ�x�S��f]}e2(S����㘙���G�l�����G��)��^K��uM5�I;��)�Bg�[+�a��(O�-�K�޼[۳;Jl�2�$����x��zY�.���#IKl'n����L�����Q��L��]�x1���r�N����k�q7|^C�Cp���\9��&�S=v�D�V.�0.;�r��v!gy����J1��\4��e���H׋�My&w]�*W�oի��3��s-�䌁�V�
���-�j�	�䩤#�W59�BP�#���o�)d�|E������G����}3D�t_�R��"�`�v�d:��$�p�p�������~"�͵&����鰬�z�z�o�.Ķ�������^eP�.
�Ut���@;�;�[�����Oq�e��
䝕�Y֛: �9 ���D��8<1{6�ų+D�CZi�%8�vG���^�v��E�٢	F������ `���#{�qxܳ����d9Vi��=H�8��q9m4b.S<r@��L?F1�]i�	A������v�eP(ਜ�4�۝%"m�s�9e-S��i,be�o��ݐ�7<VCR�쬍u�@�]�����hӡ`�9��* ��o�Ԟ�a΢����f��_��J�h�\Nq+��CS,�I�P��܎����5��]l���N�P�߮���}3d���D�Y��+�.�I؉'��觵�#��i�҈l����<���*k�a�m�*a��H̷��ȟ��hr��yf��
D�v���P��n��<"�/\�ϡů
�=R�z���(�y���b��Lf�M�4�8��n@�B:dH����\�ػ8C�
բ#��_�{�)0_0�P���Z9����F�ӭ8�Bd��|܋��kH_u�.@6�������|�`C�������M��Z��C�?�8.`'�3� ��Z�Ӯq�>�q���1w��D��v ]�JR�y���֢�7����[�X�gN��H��W���b�З�(�-pl�(���|��,>���-UQ�M�]�6=�T�k\�cny>[&ٟ���i�B�uy'�Ac���* H@�@�\D�?�ww\W�n�׏���q�l���8�-���fS���C0~�jx4:�8�Av�n�B�1��� �t����<�Κ�Ш��T��qrA���t_��^�u����W��+�C��y4�[�+[^t޿#қ���y��+����^�4*�w(ƒ��Ș1ᐦ���y+P�Ǎ�݋�(nQRn�� �R"\�]�q�. ��З�m*������K������#���8�X��$�5�ɜ��۸XY��R׽։�(5R��|�
%y�O���4k�0��j�#2��oT����f?� 2-����WER*�)�����w_]�;�D�#^�_�h���Mo=��Y��=1s"I)��j�z��V��y5��B���v�} "��a�<gʭ��&�����v.�5���G���:�nVX�R��F�z�;�{}���S���Q�WN��ʬ�6��vE꭭�$���.5���	��R���ќ+�j?~�\�c��d�R�{4n��aX{y���ĥ��%k ��!@��=8�R+�� �#+�#NDe�j����+	i%�T�h]=_X>T�a�DFѣ��*������kd>��XV��fޑ0[� [ ����d:T�`�"��ѭ��xь��| ϡj�t�}���Υ]3Z��8gm4@OV�*�aV�9ӊ)��p>[V�����
�T�0�E��J�/ʦ� �����}�*��*���.�x{���{k�n�H���h��2+��� t�Y��F���"��[�����7�����$���ʨjJ��ys���@3�ү7%w?�?��YQ�#��'��	��+W�oH��F�x����ep��{	<ݝ�	�TN�4�3�`.�,�q��{�p;LG<��=�F� �~�^�rj,N�}��.8'd5;]0渠t �$���%w�9�J��O�֗YPz?��]���ق��$��'��`L{:{ɘ�X �%)�$E��h����S�*�N������`�X��=Z��HyKG�Oi�!|Dp|�2�!�م�	�v4�֜"6�lA��u��6_�ݍ���雎J�2G\��E��l������	�8��v� �q?Ͻ9���oÏ���{�X9�F�����J��s��ͺxñ�@>�r��o����%��B�w����)[& /�\0=
fc k�g\��@V����6�RU9	��R����$m%;����y���%�f�+����"��]7�lG;U#��r���c�K�;-#������e�M�Q���O��իG�7�?F��/���A頦���W	'σ�w�;�x
A 슭ન���`�8q̌�Y�|��0�	[����y홽E.�~����mO��i�xF*q��wm���������m6��Ӊ��W������	0�%Y�yMa�5u�kb����\��!��,DM�D��~)0K�	5�u<��}����a�w��c ��M��<)���~��nY��M�rB�))O���^9�U�31��)��f�8 �<~��c���S��]osO
��e�r��J�L�9��ӟ���c�f�C�	<n/�:_2������"�����?����84�iB�ɨ!a|Hն�z��ʸ+R.�P��k@>M/Z'��a�T��lf����~�N.�lt�9���NL�8�@)�˫�2Q�d3�x�1A������\�'=Y�!��&s/���]A�_�c }.Aճft����I���V&�{��a%)�N$#�Q�����Ao���{Z�h��K�}w��������8�b�hp�.n�p�	\�+فS�NK�T���z1ѩ){Pq��# ���t
}Pڏ�T�t��`I��o"�y�ᩞ�6�Wv\Y�]P����l >����s�����G��1#Ge���T��+E�_��"�C����3n�΢|o�cL|G��Ót����A���s5�Sn�]��o�N��WрrdK#`rc��}.[8?�f�3{���܄A����2X;��_����4���t��L�٣�c��[�0D Bz����@XlxVHYEB    4f27     d40����bFx쁠�vR �3CY�D��Y��IU��AX�H4�[�^����{���K�"�韽�_ޭ�� ����-�g�Ὓ���K��=;ǋ����)�ԃ�DB��h�1��L1e�8�>G�ḥH�{Eܫ���i�H�A$��5iJH@78�@�\	����ԎC�t�l��T���e	�
�I{����kcP�Nm�_���nl[�ž���o������T��:��`�'"�E�����_��[f� �q�y�����ô�r/}1B��
����e6:�^dOk�ӊy�r����ߛ����*+�^��?���,�POm��}��:���[�G#��@<�|�3�k6�׿�:`π����j���G�� �jS����ř�y���ޱ�l8d���V7.g�8�M߫c;LL�%�*�Ԇ���[��Fi烔`�Yb�]\Si�jA�7��e<�6��k�n4#�� ���rw��+��T�����m����IO0lh|4G�E��ϬBS(Hw+2���w��_�vZ�ԭ�2�0s�'�A, �RC���ghw�h���QhyÍ��{
���v�X�骚R8K?|�~�Qg�D���l�0�x]Ҷ<_��4����5q�]LmדqYi��]�Ն�-�����߷�12�L�yR��fM� 	���nx��V��� �>�#�\T�R2�uۼu��}��S�,`Ѣ~��8c,'�N)��VfQ����<��`,��@N�ߩ,Mb�᷐���q�5�^]��V'w����^�ލ���O�c^GK���39��rA����3b����7�1#bONn�<*j�V�v�Sͭ�P3�t��P um%/sP�D��h�E�D?d!�	��aY[_��1�)$�I���
�(�)��)l��2�Y2��[���?-*ƚZx��)�@�'�0�­�;���|ZG�#����3���]$��/Zk߅�5��?�-��́��*/t��Qh)εQ�o�js)lpo�:Hv|d�ʾ��5Ca�3H����N��'n�[Rn�'�9�q������W��U���!����"�UBG�2�3�UZ�#�O����̲�ct�p�B�V�}�A�)�¬�}a3��6��.q�Q�X�jci%/Qk^�;���fh�9�g#ע/�5��6��ӷ�'CORGKV�)�����;�g�cQ15��0C��"���;-<�9x��_���A��N�Fc����7�$	��%��3��˔���}2\�x�VS���{Fs�PΣA� ��e��>Hn��atN'{M|Nq��|���x�M5A�S��!0�l+ka����$s;�d��Ĉc��0��V��L��? �^JyifNLGA��2e��o�����洃��p�X��
���<([��xQm�5S:���a��Q��?�)(}T�LQ~q�qZӈzՂ�Re�,�����kM��4l�.I�y[�K��4!~ϟ�ւ��촻e`?�7�������n��-k�k8ģ����bX��!�Rr�No藝�ZO�9!΍*�����:�d>(ԋ3pxÀ��pk��1��9u_�عY��N0k�7�X������o��Ҕ(�s�r
�s���X�]��Eg)MiV.-EW���	��O��m$�G ��
�OV�w4��H0=o{?��;�����p��Nuk-��c|��綔i̽��Y�Z�ͣ��{	)�cD�ܛu!�Π&C�$gMA��ݷ��Ǽ���`���|T3,���%��8�pz��}$K��]�s#*&��â�C�vx��v̆l�g�z�dY):�1@��;'͏z��H~�ꁿ���ƴ��@�,}tS�.��DQ�9�c������c��˳��"V��9�������_stJ8X��5C4����A}�q�Z��x����.�fC+y������vB%�]�1_M���פ��D�64U���Ja?K�=NLn���A |��t*k��~5^1�]Έ�o35Q��"��~q�|��䒞`ꈐ%�J���c
��eh�S)��(^�Y:��뛷����k����d{'NW�5-�)B9q�[���c������P�b�X��72  �E���="{Օ<j?L�!�8�@��:��Z���i7�E=�6�8��[HX,Y��"�1ͧ���᜹ �ǹ26�ձ{0�g��s�6���w9G�Z%
 �W�M�N�3�,�Y4J�|�?bdQ�=.��kw�;����н���m�OH��&�:?�9f�
x����1*CO���2n��K�� ���X��9�GKIx
VEˏ�/e2V�7��/e hv6X��3"��lb>��ɕ���LPą�a�䪃�t炙@�����J;��v�z��g�ݺoAK
�1ao�QD�<Ё��n��Ҳ,k[y0�Ny5��	�n�l�%�>Kxy��#��L�2�]au,B�1�;�$���[�ZN����(�:puy7Mv��D���=�yq{T&tpk������_L��O��~lX�+;�������΢�����$��]������6(Bc�����������"v�"�{̄���F=C���Y
[�g�����Q M)7�9�+s�$mM� �K�SnĬ���3 �=�7�!,H�_�|[� ������*h[y��Rr��2�T@���ڗ��N��s�=jG�]�	q0[��U۶e�r�P��!B��*Xh�!2�_Hx��� ����}�X7 PTUh���d��ӷw<�I5��F}_i�(����E�d ��n�IF�`��;h��=�W�b&�0wm����5��4�*�Bf~�4��v؛2ǇY��H(_�k��N+�:�K�2��.h��vp/���Gw�Q����P�;-�)�Lϒ���{d�ܶ)C��! Eq�I���R��_� ����8�۾����
l_�h���1}5�up��a~�?FP������Ac9}�{
n =��8�M{��
	��F�4�jG���Q� \���T;�M��[.��X�Rq�+�L�u{;5���I��J���Z�nL�<m~" �K�Q�P�0��IdPy�=����e��\��o�/���뉳�{�y���j��1�(�\�j[�;rܝ���Kd�hUz���	��8�aj�<iOueS�=����</:!�	�xЛ���}{��~�:�`H��~ȔN��xp@�a��,��
=��H��b�z�䶹R�M�Qi'�"%����и�@�&>004�+��)�@O�l�SnFy�^�bM��Xbϩ�W�Ҧ*�0g��d9�r��ް	訴��P����7�����-�Ul+�/�T<���3�D��綺'�&�-�tS�"j�cc6�tY�|���%