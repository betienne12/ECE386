XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�]a��n3@��%�AT�VuH���=�}�2lv���~_��7#�.�q��s�uZ� 5�l��i[��#����82B�H��HhE�j�6��ZE�'�j�9�	���#����q����}�B�eȬ|[Ǿ�]�rN��N& MP��/�� �R�(3,��I�MOW��2��P���Mָ�~��]%yt
O8�/E,���z)B��}2��ک~3�J�&����J���[�C|���mE���![O+�v���'�� ]d�p�_n�P� d���!OO�֧׏�0e�Gh�^�sU�����* �L�����>��Ɠp�:T��s�{�X����'+f�۫2y�ʨ��.<�4�~���)��ݞ[&Q�օ�A�#P)�&7p������k�'f�h�φ'����f]��PVd��G3q���$���r��`Y(�S;��^;}��>�	{ϣw�Fs���l��&�-N��]�Bd�1/�-`��v�����2�2� stvS��%���
���c�{F��~�B����^�W_J{ycC-���Y�oDdM�<}s�F��0�q�J�#�7��סo=`���d������.py��2�&��'KNK��@�}�徧�M1�sn��KK�s򽚜W�7Dm[�ܦ�����Ļ�����.,̃t��CNĉ�V�ލ֋�Zk���4�ƺPfd���Ml|,46�XUgP�@�O����3�F�L���[	%_�i<�#�%�e�:��O�߶A���� �"F�J�܌9��!��ϹMXlxVHYEB    fa00    2480�Wj��5fGC��8Y-7M��/t��JK]0W �ii|/?�Qv�N�.�eU�s� 3A�m��Z`u[/��]P���O�	�Y��+zj6�0>>$8i��2W�T&KmF�o�oC�(YKH?�W�N�ϣE��ަIm� .<R\yX)==�]Δ����=L��$��+�Q�M�m�V!�҄v���vg�
�������� ��O�Fhs�)�~gS(l��ɝ4K4����(<��\dv�6�o��e�Je� ��koCt�P���:�Rk��{����ݍρ���W��G����1��$n���M�~9���T���5$��uA
gb�G�a6���`��I��vS˞�9b�
*?�Rռ}m�5sB���%w����EN����j-�;$�g9_� ����O\h1yd�=|�	L������ #Z�eߙEx�6a���S)�L���5r��96�
����v���\�/�n�^6Y��h0��3�U�4D@M���t"9�4�ӿr]:9z��2���� �.붫�BY���@^4k����Ǥ��`Km<�J;=�����\�!W�Hd�]0���4�b?^1����@f{:������}mֻ��Lḋ*��xۺ�8��Fq')C9`���$o�	��@}�z�O����]����5l��H�ź�8B�-"H�$���u���җG��_/��*}0@����/WQ8ꞧS��UA�k����u7�q�yϷ}���0�F�6bh4���:\s��h؎R'��~��:���Ǳ)����t�4w��#r���y
~�֓b>��`�i�9�O����T� ��g������l�ߏ�m�����/���Nx�f����MN�Vٲ�iW�ڲ��r��׊?��CKQ'�E̠���,�;�p�\���l�,��-Zs��y�ip�o�U)M]�O��&�G)�ȑ��XO.��AL�*3���vN /�x��r:͕��ӝ�5���TI=�+��zAg�^�S��B㤙�P�#Mm�@_� >~��3����p۫εr�ƶ�Xz��T�F>.f38���,)�[f[ZB����|���=������;�4n�@V��տ�|Z��adq��t�%�����~ִ��4n¬�jA3�,��c�;��	��ڳ��J��?A�A�|�Z�`1"B�K_���Z�6i��c�^-��0*��3,����W����ۨ��gW��~;U�ď+�ep��SA*�n�E�ݹc��˼!�y�p|��m�����$ʟ�3J��LOO7��t��:��>�JAf���p��/^�5��K H�vzH�{�ܾeŅW_Ŋ/M@�!�`�2�s���i��'NH���[?,B�ח�tA�3*�M_�Hљ?��(*��a�ځ�`vO=���[c�l�L���g�i��Rd��5Jufb<_��8�L��%_j�k�C���p�D�o��Ȟq̦��e���]<M~�R�紘��I�"k��c��Ǚd�N5��a�%�0�Q]2���x��	 ��3�B��GK���@D7�����K��m �/�볒[v��]
�F��x��o"T��}nF�B���/��յ�S�^�&#[�E�^F������u]�G��~��8$�Û��O؋�w�U�D��ua��x45��+9U�`�v��g
e�v�2�;An���8��ب�@r^����oS��2<��O�f)�B��0���N^J�i�.�|���p[û��"X
��#�B�,m\�c�bjOD��ᾢ��3�Qp���g��1,������^hJCLی�G%0�/_���f}����a��E���S�R�t���G
�������\9�4�d�h����x�R)�l}�k�|��ҧ���ZV������T�Tܚ��.�q((xk��k/�eE$e4�	��5� ��ÝF4_S&-�zY4���z���;S�_��>�E��F��}������Y쑇
�1������m6�������x�,�=�ǰ5��S��$�%Za��
�x�X��&F�l��X�i+F�F�ki��6�*+���}pUM��:|]81�"NF8ݑI����k�^����.a�&$�,K�}���h1�[z�/��|Q�TSɛ;C�7�w���8v�
�>7�.;��U���YHp��\�t0	��:t�j+���b�ư�yVڛ�Q&�D�%������u�y����w�F��wBZ�NF��b�~�?6�l�f�Q|%��`�l5|uՌ�޶1N�ӧL�ʥ�J�`���Զ#��S�zh�
�����6�m;�Gߘ��|�1��E��`������Ж_�$-����d)K�hS~H��`��e�^G�Ǟ�\݅-]@�
�*]��Z5"@���@bX({ND������@)O�%H�#}�С��~���ˢJ])<�� ���a��g��b�+%�����`���f��B�^�*@b��Ac��o��o��\��O+�%' W��@��e�FC�~��u���g�u��𘵊 ੿�,և�ic�����}8�H�h�|���p.��j�$sH�
���!�Ɇ�K�a�U��*[6kf�j��hb�|N�À9ei�uUO:�n�\nT��W�x/d���mE� �2�	��+� �b�������ag!���r�Ez���b�̳U�@�"�{�=s��1H'{\�'1\�m$�jG��y����nc��e�b":�qG?8��uU3T��z;�	ط���@���@�R��l�!L/*�lU�!����;�E3\^kS����ꌽ�OISܯH��֔�m1� w��OX������O����8�L!߄�������Y����-�PU�|���uT�8e]ߍ{]�J�����xw3�ɑ}�צ:��v^C3]����5�K��\�:��n8J�:y�D������y��:b���5����S"�ר�圳��~d��἟�)z�:�� � �n
(J���;n�<^�\s�^{��ġ6(�#���-��7ԣ[N�f'���*%�u�JلR� ��/�qe���m�M���J�+�]���Xx�SQ�mQ�yi���Z�px��r-������,�IB��;r:��ҹU�Ѱ�z��)����&95�훣�^�QL��^��G MtO�>�PWQ��Ѥ��(% o\LY��*u-ٽ��!��G:�c��{�hKf`J�Z�
qz���p��rjt�3�w~Ы��,��*p�Ҹá��gڝ8���89�CK�ht��-�,�LN��[}/��Oa[9W��)�'���v�m�̪ndr���z����2�W>�lͱq4�֙�j�[����V):��|:�U��X-#8���麫���1N�Pjߡ23�}�����B=_!��jͣH�z�-l��[��s�ꑁ 
�wm�{NL���Ԟ�;�V�P@�:x]=Z�`��	�u������Ò�7kw&˃HHM hO{��o����i!��x�����9Ir-���uyO�ٝ���w�L��)��^V�ޯ���ya���ߦ%�x�t��c{����f���9,� �����Mp���HL@8)Z3^�m�H��0��b<���֏n�dR��g���"���H�:|P���iL%�wE8�-"��R���_�E�^�<2y�2�K��Z�t�>1����x��5p+��{ G+G*S�҅�`��e��
��u,�i�#�hl�r���x�(���] Ġ�sY!w�?�nؑ2��o�o�'�'��.�oM��gb�D������N���0ac�/�;,:�E3P��ü�T��g�b���Z>t�En��կ�x\|r�$�zpa��B��xʯJ��FޞCL!vA�y%���JS����&Ҟ_Y9ț�q;06��c�)I���U\W�&�ZJ�vyh�bA�(�`0� (���;M��',�����ͼѕu��ꝨZ� �)�%�H&��j$���0ɻ��!wZ�n>�� k�S�C̴"G,X�ON����▵5v&��~bӥ"�];00J'����O ��I��O�d)��� d՘#C��ٺ�(����(�j����b���|�מ��r3�KX�NDӠ�(��?O�%~`�����&�_ �Uw!Mg���U����W���_%cl����ω�)��0��^���/�(�(ZW"(���x&���'JC��q@Q�Mv��g�4��|��o�AF��KCJ���gQ$R����f"r��8����z���?NL�TA�W!Gd��7�}���V�Vs�k�B��a۲�׮�Xl�Lûi�����r��͙�+�'��P�j������#���9r��'U�i�eD�́PX |�g�F_ӵh��o�~z\@Yڳc�&��*7Nf�i��T�D`���^����Hh	)�u3,-��Zڽn���p��[�����m�������.���7��k��^���z.VR0��m����h4(i�6�%Җ�c�}��s��cl3?N��ԕ LV����dg�~ZV������)�*�msb��b�x/?��߷pl�
�f�5] sc�:"���-�8��aܡ4�U���6B����آ8F���uK�r���j��-�>`����g&�y�����_!�� 5]�v�en�D:�"ܓ�<�T�!���`��vh �)��D�\g�*`
�K���Cڢ�3ꖙ��,�X�i$�m��]\a'f� A���׌��%���cB�4�Kpx�X�é�%�Q ��E.#��[?�>f��Y��B�'׻�F��S@гJ̢
������hҿ�BN�*�-��߃T�-��U�)�v��-����*��v��v	��=H$.�:�䤨g)v<ðY8��i��㪍��/��d\���yM��B��8Mk &�F�����=�Q�7��F��y3� ��1︧���pu��.'�E�|.9�l�	��}���o-A*A�L�������l���ݍǯ�Ⰿ^g�<�6�r���@h+W�GQ9=N�J0�\���k�)���o��sV��i�DxS��3zl���� ԁ�*�^�1�����) <�<q�zzo�aL�?�9��g��ftP�,���:��(�"�./c�i��5�ak�~��˘��	!�6=3�B,|5.�q�]�o�?����Ȃg�|K�6Y�{TW�����K�*��R��Y�G0�lw��cO 8ӫ�+�H׵]����˷Uc� ��d��`�`���9o���W��u�2QY�L)�����I���N�p
��k�%��`�C������V��S��%�-G/�q!�j��O��duv�sb�f:����NV�hc�84ВB���kn�	����Q��c1���_KK�d�����j		WP��x0E�xO�t*��U�V#��W#Z_VE~��.R��YE�'>c��љ�f$K�"������~Gw��}�:I)���W�P�K�~!!��K6�X�����V��m�Gb'�;l������"\MI�.�+e�&"� �i�*���q>do�Z]r�����kJ�"�� %��9�z�_ �I	F�+EܷN��t|��x?�:������jFCC'���j�U�(+�y���t��Z�ڈ3Bo�*8�vJ��o�n9�y��@�d�:7�cO�#H����
$BR˟�8��/�9�0i0�"��Q��]"�h߻�jS����E���Ϣ��ȵ���L�vw����OfC7JM�]Afӫ}�;j��O\��oLYO�m&=��!"~�_,o(� ӫ^��>��V,!/ͨ���9��n�4H�
U0oD�#�9��
`��!�˃������u§Ţ�Qx~�d@�GO�Sgҕ��;ߨ`�@�T����f�kG�.qC���B�l�ij�����*�-����`��`#Ylp,�_|fGG��S�������P�4$���,<rO���
,{��k� 鍛������朰�okm>��-�)���q󯁜|��4Z����Fl�UrL���-�5�2y�L��a=��)&WT�͚���=����ز��]�0���v5t��5��u5QP�</sR�ޔ�����*����+7x�=d�`!��(S��X,�f�w��YA�N���ul�Vν���]���e�0F3��#�-j���,˯���x� u�M�,9Ղ׈�n��2͗k?h�R)�%�'����K��p�z�f���!��K�$� ���6_�cx3�/���4�"o�*
:�����лcCu�Q��'�k�كQČ�?퀢9cq�ލ�������¤ͳV9��%�<���W�I�Ί1x�Āp����V��+�f�i�hZ^�������u���1�����7�#�k*��rw�$�/�9Q�'�����ˡ�~ɜ�
�B�=����z�Mh7�P�F��l��+'��yEP(}Vڹ�_�^��E��w��hW8?�KA8}�	�(֫A����IU�^���Ë�T��O"}�8�O�2�@X�vF�0�8b���2���y��t� o9s]���9!�lzˣZ"�p��lM��n"��I���Z�=��go��}�WԄ����J�V�[�ej�b�p��-߉2QȓԱS ��t�钰����	��x�lX�s�v�O�@$�;	��;��qA�ܮkoPN�MY��<���s�Y���
�O<`�>P�E�������wY�~��d3�Ց�1��P�D촳�������-�s>�2�αt]�n�(�C���'�,������PӨ$���2+��(���gv���!�i�~�+�j�@.�6Bk���"d�J�\��ջKx�&�L�?U��_@��^0��e����֝�Gә����s,�����W!��L<[���5Y4Q�����x��k*R��0��K�
n<���E�=(���}IO��þ<�%A��A�������a����S~��@�DQvy�H=N�D4^D�QUFw�'���~���^��g����rW|��ӽaվȳ�ޝ�su`0���4�"S`�0�K�o�ȹ0�K�� :�|�U'Q`�]��FL�a�D�u^cw�^kf=��ٳ�W�r�4+v����ѧ~v�"�2Ь�N)HQ5�f��B�7�� �{N|��a�C	�# �!�"�����g�H��G���V)`�"�g9��:��T��^p`�nz'�d,�$eaq�6����.���ʝ^�#�>�,,�y]1�Z����i���:wˏ�Pc�`ǧ�{�� !�09+�Q�hYrG�k�Q���l�Nif#R%p���&71���&�H�@�UMf%ʈ������5Z�HS���=k��}(���GrL'p�7��4��'~�4�H�x5��T%ygdנ�~�~F����4��T�1�8Q�g,ʭ8a��?��Q_�.
"���"�ʂޙ� 	͖��b.�=����9y3z8#�޸6k1.qiw`Aݝ��_!��a	�%(nWh���y������O��+QýߑØ�3�4k서وz��.7K��v�G_�K� ��ll"ܯl�]��/���8	w��VqU`���4?����F˩��"����	IK�m�z�@��^6*2���E4B�b�6�ת�o��T���w��tݱ�	u4#�*?�[�:�	�6�=u����wz�5�F���\P�P+�V>��{t��πL�����p}�@X�=��YF�C���27���T2a:��a�'_��$%.��T>��8A`Ō�v4W@l�NUm{���z�R�$ ��� �^G�?z�O�`�##yrMt�޵4��N���ScF7Ry�Yq�Z�O�A���.��?,R�ǃt:�3�k�&���`%��|�MV��S��?`(���R��`!�^����p�� ��8*=޽��A�w�K^#�/	�f�2'�9V������
�<Ж�6ZK7��̈�\E(� ��P�E�B�ҪYu�=O��!����p�K.H��M�`D�,�Kb*���#�� �4x8ŭb^y���������K��W�)X:.�k`dcW�#}q�����ݴ�����
]�XU`Q*�-������ ;�b��\���d��)��{���j~��1[I�N�{c쥵&J&�S��6�gV���2�LeK$$=����JV&��w��Zd��5F�ҭ���M��v�9�.L�A1PWuD��f3FK�`}�B�	�^U���A�I�4:��^���ڲ�D'(oD]�>_���zwY�X�T�'����_�;P:T=�ծ&�¦�v;�"�y<~��'�nk��=��~��{Q�6��-s�a�n�x�<JrꜲ���tb�0w��S��(ЬP��1��u[Ј��z�"��B�Vu�慈��h�m�����a~�9?�z�}V��$�o =�b���}���Sd7<�\	�g���C/���!}����Q�-�z�z���ڤ���g�-����{G�#��e��L�+�?&V�K�ś���۝���$d��̈��A.��i�b#�D�q��l�>I"���|���Y@�(]l��QǼ���n���d�\�Z�T��K�-��k?��8-�
�oԜ�3TY��s�;��좟hp/L��;��G�&��Nm�*K�n7E�k��U��B>��Q���Z逞GmF��ʊ �@'��B�̈́��f���~z	Ue,�Xl<|��`?��+L|��!���4�0<�pL���� �]k�g�\�/�2J�ߙڣCXTE��Zk^'��(��|3��b�
8��N"���8��$�C5�B034J�̀"��W��$�9a�;4M!@��Пyg�������)1%�!�B�]���Ra�|�j�1!gO�g2|j��M��Ѓ�X���d�R��xnĵ�;1W���[j��,�b8�,ªY9T�� ��Z��,gH����f�~���6wma�sN���/q.RJm?={}� 0M�/>�i��\�&�}'�Z%0!I�r~�¹t)���C$wl�:�g?A�]��
�{H����s��י��M��>Z+�}� Y-�oԬKJqjS.5
;����6�H.xe68Tl��8l(��]k
���v	<��F��
���6�m�.V�Z�;q*_߳�SS(�^����Kve��pܴ�b�e�p<�������@�&��}��5�F"Hi�W���Ƕ�� �nu����m.�$R���g<�C	~Zх�e�h�F$��U��7�V�»>���=5ài+UJ��6��{g�%,�+<Y�)���`X-��mT��(_���>���YWZP���i�2;��/���
dθQ�XlxVHYEB    964e    1150"�����jZ{����pT�N�^A;\�47�dc�J��!�.�!�cB�i�π8����^��s��v�4�ӻv��Q��	Kj�9d�PBj�s���">�Qص ��%x=�D"�ܜ��v�n#�Ӆ�&�y�<"��\@�8�{���P���
DO�2�nU0F�y�.���j�N��Deot�Wmd�oF����ή(Nrt�&�W���r�ؔ`\v!����G=J_�4E�'����>�Ka�xuH��
V[r�b���1���g��#IځN������Cl�j�L�W���!+ 2�SM�5�%�m����J�dIcL���4����z����C��F���}�6rh������-|>�/&�-��[�l��˅� ���4�*�y�\>��n���Ě�1�xu�=9d���t"*��_�~��dk�x>�!�˳Z8q~.+wnl�!��u^1��'��j~�z9خ$L"���� ��|���_��o���iTL�4�<�a��^� ��)#<��TFs��,��}��y4�L�B�k��\R��o�?�*�-Ƕ��(r+Qw�Kͬ���4�?5g��F�M��x�#�%{�����9�~���A�A��)�:.�N�{`���}
�ѫ59��$8H�&���r��ǋ�o�Ɏ@!���k��(����7�D��c6��|ȟ1uJ�WX�!�%�Y��_�� �����}U��O�O	���¤턊�2�Y>���)�J�d`i2R洏�%k�K��z�����=r3����]���e��Ql'�c�>�4��F_>����q�۾�_�3�v��&w���#�#7>|�@����m�gW;VP쏍��e�ڀh�`���S��'�FX]CtT����xb�t�-�^�{z�J{�k~�T�ҲOˉOL��2�*�~��!dQ��G�I1p�^�[�Ɵ,'��]%ł�U�^��j�}�(�	%|H���}�r����(����Ǒ+CU�f�Tsͤe'�>���ư��6��չ3��A�(�X�R�&��L��8��XV�zf����@˪3wS�� )#��?�zt�럱�]0�>͓�3��n�)΀�d���Òv�iM(h��!�/ľ��������l���>��C�1-e�Q#=�p�y�j�̸W�[��)�|��!`��������A�i�֬�h�J����@���F;	�ay�o��.J�.
���<�0B��f�W�����m��
��>Y�k�:����j�voo�c���ܡ����|= ����#��Ʌ_�cb��b���͜M�ɦ0��cFCZs�'�ȅ�#l7S�7E@G�n����!���<5���ۻ��u{��ߟ�E}ɰ��;���8�,�p�slqg�Iyl�ge��}������� �G8M/��M ��NvZ���}F}v�]�?�ݬl���G���7��l�r��t���T�;~��L�~�[¾�j��o4��W��r��"�W�zn|�k��d���+b��_�gi����_z�c-+�h�bW�yF� �]�?{z䉧�����&' ��vVV�Օ��0M���$5Hh2X���@����U���q��1^�30 | (�V����݆��ij8�;���t��K�uEu�F|`D��-����P�ӉB`�]t` � g�B\T��'��?f:�H�lʘ�gD��|��	�:V�c��w�=ǢY��)���H�$��D��J�/"{$�Zb�(P���A:Ue	�v��2|�Ҿv�f�ɤL:-F��)/b'��8<xѴ1v��E�<@�Q�mo�o�6�ܩ3[�m�YV��z
˕vpC�v�f�C�����I��T`�(j*�ƥWjBdA���O��~�vL07&&��>S�F� c�|�-'C�u��>��[��;�EK� <��	ɓ)�
���']�?HT��
��*6�.���Sx&Л����cR��بp��9Edo4�rс�*��x��N.C��K��.?������&����zep���<�����_RX�P��(2��1�4�v=d��+�8�F�7�wPt��n����K4���;
�!`�C�zT��D�EȒ ���q ����/���@�vd�1$��.�5\��V*����m�[j�+'T������^	_�S	�/��i�"����.[��m`�7T�tz^���EN g�]�� �W6^���>�1"���Og+�ɳQ�vG4���1���ўǻ/rу����#��X>,m�N�~����Gi�0
x-��f�����l��M�)��B=�R�u�ͳ��\[7o�l�]��Eќ=l�Nsw�2;?|����BH�e�q�s�T;���7��a�\ʙ��x�����T�<[�\�f����V�]�o4�8�</�0q؉�2�RQ*{~H�\Y�Nlt�M�R�'WN�<��Jo���Akp&c>h���P�}s��!�a��0��c���l�h�=�S�|�v���V����Q���+�y�o���7����x'�:��2�A�K�Vb���P~��<��OYy�rؔ�{	����"���%ݿl�/zh��R�f+�0���6������ѥ2�&��/�J�}��g���{7Xn�c���.�Ӿ�"�w:����
�8XQ�wC1������H�(�	�������4ay�k}D����B��'��>w:a!f.FĄ��mW������1�<d{�vp�	ly2 Cs�W<�5��r�F�d����sȴ]�hU�C9S��I�X!�h֞��L��#/@
�=)z�|����s��8C{Pa��83ũS����1�ҫ��y�����j/�<=�/�tK�Hs��w�����藲=fm�[�~P��쯰�¢+��%1���R��+Cz"�-�[(�F,s[w��T_B�%�V{`4���jE�A��&4���g6.�!���ZȌ-ں��䝛�����Kvk�5σ���c�r=�w�R�߃��	rޚ8j�)�8����v��ŏy����N���*]b`;;T�M�7�R�Ҋ�M<�9��z����o�|���$���Šwn��H���*�X�W����H��V���#n�\�U'K�Dl�����3�A�)�mieGQ�&E'�
æ�K�����
NXvC.(��s��u����8񱬹��#Cw
�%���zk��Q����I�^+"N����s-�$�S2D�l9Μ���'�����MC�G{�L(�E�q�R��D.+ʁ���N�R�UM��]��]ꫜCz��8����5w�7U=t�"p){���'�.��;�Y�y_ L��_Ч�![y�m��)�8��b�e����j4�1!oHm�B�ѯGV=��5��i~�l����jx����8�ԓ��g�Ч��Q����cl�-f$#ۯdc��T�r�8.^�S-�9��ա��]��S������O����^l���!5�Wj��o$�@��f��`A����+�~�rg�c�|*%;���ܵ"y<O����g[u� �	.$m~�|�y��Jo��D�f+&�Od�υ��^U�ȶ� ��?3��qj��I"��R��C��ɡ�_��(r�P�NL�<�A	��²+�3W���P��n9�}@�C�=��w�	��g�J<-:�D�V/0�4�l��U��/bz�XEM��k���Px~�����=ҩ���e��0�WA�3B���I���4�̌O|��L-��u	�Q�[�����(�,�OY����-
x��؞W(�~��M(s���l}u��Ҡ�e�Td�u&rx��gO�}�}T[�lj�0 �eX!i璑�|�M pP�7�#�U��*[اfC�����ԊU8�e�eC�|�t�j!���$5~C�g���:�Djg�:��{OU�v��]] c�Ge��.�H�~�������g��E����_�@�!�k^��ެ�XF7�B�z��9aH:Q/+�{�BR*ݠh�]=�D�g/`�g�X�o8yY���,�\r �zgtӍ��nm/�a�|��l5/��qc��9M�}A��ܾ���������+&��L�(����e��g:�-ȧ�b��m�_xd?7�30X�C�6n�H�T�N�t��7z�x'�;��A
��u�VkĂ�hR||��@f��s��.g�ۚ'���|�[b�C�O'O���pʄf��;��o�-P��Lq�d�,�u�,�mM���R���?��P���\��DzfԈ8�����3f�Ƈ�ͻ��_�9�j�v|����#����q�.���6Es��&E��h�r#c;$cS���z�Q��Q���.�����zg�(
#Y��_�y�d��!2&G{VH��N�? �$$N��&��^F�f�0+`y,��xv����Ue������