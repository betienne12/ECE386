XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l���c0K��8τx�=���!�Z�i,�-}�T�!3�(����b1eb�BL��eo��P�am�����hR�[���v�PC{sn����$���)��ɞT���"������=o
�>��՗DKw{%	���i:	�nѾ��VS9'�~¦���Q���a�O��F��*��H��!�=�	O�����{�G�4�ІR<����t��$���]C���ٞ����=fw��N��)����S��ʗH4��w��-�u�tgD�������b8Q�%�l@����������
\_�x�������@�ݝ�Nfh٘P���상�켉r����m��̈c�hN-��j���=����¯ġ"�n���\���6W���S#�� jn<���u�:@��#����^��𼶉P�6����+�HUbS�l�cČ�0��1-2qQZR՝2B���hU�bݡZ\��#��ң�2�S�c�Sd-f��2Tq��I[]�+Qig)� �Uc}[�e��}��7Q�eu�u�|n�sx�Ǘ��~؏����*�SDw+��j*0�c}�FDWυ���ap�-�*�G�p����;Y�I>B���|]2�.{W��,��Kmݼ��?;-qh����`�~�R���4��Å��i���-�9�hZX����sRY�,d��v���r���4�%!: �,�QNZ`�pZ���9?8Y_� (qz�J�p��B&�T�O�$�D�c��V$�5���_�	�##i�Ӷ���e��XlxVHYEB    29da     af0�0�� P:쫹(���x�/�i�G`ZS��6rMƳ-�_w��m�n���V�-_!'�)b\��v�@:���: HOy2H�E���(�.F�W�	Vy=��n��^��x;�ⓗ�t��מ8��]Ѕ�ev�E~o��K6k����%ߐ��	�� fh������V˱��2�m��E�t�i��j4��j��k̏��9�4���Jk���N\Yu� ��џ܇v�S�5����:�D 8/+���T-Uh�]�f�Ѻh��f�2�j��N;�"�Q���h�Pej��l{m�S%�T��`��"s�Eq�ʔv:�jyP+�u�\�l�-�D�P�w�15�@/38�	�z� �KR��C��;}U&��'�$��̈j�HtF��;Wf�R�O�,���c��d��r�p�_��U$�KC�Q(밑��Fcu�/h�Q��2��Pm�iV�u_�����ג}��p^���5� ogm����8��w���O�E[���Ɛf`��,f�bc�Ɓ����N�,K��\��w�@{��<ʲ\y�i
���(a���H��ɏ��K>5H)/��2����Y*�m;�w�:�����<ićb�RmR�YX�U�7�J�kY�^7x��q�,M�n�r3t�-�Љv%a_h�IgÑ���@�8�*�et0gJ�p��8�4逌��<�U�}��(~��MM<�?4�$�Q���A�,g�|��M����	JN�A���/�)��<u@
wi>���g��+X�>���Y��&؞�h|n�#�FԿi�3�?�����F� P�9�e�\nJ#�7��C��X��x��b'ʮ��D ق�) �i�������cM�A��
e	S�M�M�t����Q�HL�#�[1Ov^���0��>��/c�F�#�+��shc��`i�}e�C�C</H�0Cǳz�+�Y��S���B�0��-��툖�!����{y��b�,�E��i
|i�*�(	����hOoF�S�� ��M��_@6-t���OgrBgt"�^ۙ%�z�R#w��t� һ�-���{6�rȦ?#l�-���;��>�=�4��v�?҄`i�qi>��������D�X	���B��G		nN���0��P$�&3|N���H���B�;���E�kל�?݈�J��x�q*Ve����ܤ-`�e����ں\�$�B��m9����QZ��ޕ������z<���qaOd��1/��s��F���̦�$��p�6L7�Z���)ۗ-�@��@�?�OS�(�՜���ʴ.��V��"�ƚnC��������h�b�l�c��������f��{�LD��DI���Hz~�͆1m�D͙-V�3M�Cmm�OS��$��k��Z�kH}�T�/j������Z^�~��mĠ0���}�h��Z�KĂZ�v_68~I�H�
�pN�@W�C|��� �@�5�	41�ܒ��j��o���1I���1�-B� ����~�@xN��U���h�fs�srn��]�����o��)��Yg��-������ܽ[�j�R�(�d�b��P _"���U��?������UV0��m��]�Q*� :E�<�����&,�]�1M��\��ά�p�C[l�-L��!��ܽnٟ 
�*ؾ��Q��L�-�W��`D�<Cf��f���[yWk�����۩fE��p�D䃝O�5�8E(K�S��S��{�Z\W[�O~*�؞�QjU�?V�������߰���n��!��l[��	4�Bh�>}��uuK����o��U�󂬞�m�!�� ��5�j�� h�'�����?~���֐B��dO(E�}l<�!uQ�Z+�t��g\���] y��J�	$\h�?w�-|k�$�b�zOy}�3
*�aMz���=m��}J������@�80ъ8x�X4�WȀ��o2E2|堨���>2�	z�yi��/�����rU�x�����w#ù��|w���uB��y�Z�0N�e����Q�?�\�� ?�|�X�e��R72'�k�*�A���h��zFwZ\2r~��ٺݏ���p��;��֬��(�ϛ^5F��$71?��͇+\��,o|�̧�i��|���(���3d��~����gԥ��B��		���Q������D�o�ĝ<�q��S:��߸��_D��=�Z�]	���?���
����M��;-�Y�n��Ͷ}�Y�Nq��ט^���Yz����57e�-0��`��2H�&�Sy��>�+m�q&9�u�I֍�|��2ob���M"k��t��\���f+5�pv��aq��F��1�m7!����;���[�K�b��(2 $�?�K̍^q�:��4]a��N(e�0�r�@fh�R� 濝���'���N�	�]�-`N��ZS�����o�KB�Qe�K>��Md�F���I�.	D�q��"J)��mM"�.V@�,�����[�.��Z>�����!�~�O�/�$��#ĕ�b�?Sj*�5��b]lv��Bc���������H;n2ݤWnf�9G�b��8M��p`�H8��.y�#��c�Q�V�qU�c��-_�|����o��}��Y��f��F����/?�V>���X�~��=��&��Y��up�'F���ל���zyг;4�)���O&�1J�~ѡ�FᏎ� n��1"�QY/�i�w�`�k�ީVP���L��rG�