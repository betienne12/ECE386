XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;��Z�l������dֻâ�!��;�3}�:�UXP�D�������4��� �Ï&��D��W�jN�u���䥐�������q>�/h�6�0�1˵�t�w�����za[d�8��Tg'M��D��y,�Dj�nXd�t���*��>���Ͷ���0V�`Ĕ�z����혌f5;��e�)���D��MI��+2�]�\3p��X���re��?랐ׇ��������{tbFn��p����0l�ns$��0Q��<�_:+=#��4R�"�A���з�T>M������"�a�#ŕ����*܊2�`s�-H�����tH��?�v;�1�w�7�Ǔ(����;xս�	��y�t�I:.39՜f�~�_/��`N ��,�\��rN��mcXS�R����U�-. +��[�R�p=��w��q�DKCS��j��5����V���sk�c����N�j��p��O�≔1����&iv����?Xn��Eyw6��u����r񑧍�u����6���0w^�Y�p_�(XO�QC���5%��
H�$���O�s-��o5<~�pi]>oL^���U#����iU�>��tΈ������Wޜ��u����eʼ�h�W���T�/A�d�x��c�fj{A�g�@<mV������pv͡�����b#���B"Y�%�-�Gn��@�o*õ���O<#��r2j�2��7`�ᵂI��'	 ��cnCo�^�e��n�C�\��v2�6��xH��?t�9�XlxVHYEB    b631    1a00e�"P���F21+��N�JzQ�N �>SE�)�\�?��wJh������G�d�{<>�68
(�ﱚ��L0�_^������G�3����0� V)�P"k{��	�VV���u�,�NN��z&�L�{��#S\�R@�STt���`YCvB�'E�K�FL���b.���������Jz�m(`X�c!@Ù<�3�Ȼ����7y ���<aa�w�V˶R<�N� MU��tP�5F�{e�������a�l#��f���!��)W�Qk�&��5�N�t�bi�xB�Nv�=����?{�ݘ�{A9$�û��h¿��c#��B�G�>���S�6l�9R'ńa�LŐe;q�7�Y�^�Z��pIQ�w��S�|$���g� X���;g]6�~?;��O)�I�������#��'x�%e)x�Y��/�W�;>*���[0���JI�#(��S��zx�-ÑiV],���b����e��b�O�iD'^g�i1�E��J�Hl��6���]��K0Ze����\���-#7S�����&߫d^��jv��~k	_�����a����#�����	�.�����#���Խ+��%^��qa���')>~��l�l�$��k�����~n��ud���?�i��pF�z%b(S$�}��cT�;�Ɍt{��.�3f.e�Ru@�2�L���O��&�6�MHC�"�Z��A���V]ζ�sG�mK�$���VT�Tt9�]�b��nD�K@J�c4M�!.�O�gޘ��>���RR?�W��.r�y�!�BL����NZШ�9\5�����]�+��r��"��!U�ྫDb�� !:���DJH&��7Ը
&���Yb���Kx+L}E��:��I���M�P�}����e���~C���a�s�����ڔ��@b�{{}F�]��YY�KX�?.�I�#B]�5�Q`���ࣄ��؏�Lڥ�ڙ�kݽ
�B�$��}�q~a��0��W?c@�`�p|�F�Z�i��q��J=h'�m^'Q���c�gC[i"p�}�4��8�K��Ͱ�]Qt�������}7���ɫ�:�F�X�h&�D�d`r��*f���8��h��H2�G�= � k�\l@��:sS[����b�)1lS#1]���W��o����^
2���T���/�����9�������x���dD��'����#q�B��^;v�E��b�g6oT��� ��{E�?"	�xؘ7�{�!A��4G�φ�d|���x 	Ϛ|�k�0dWفP>W���>��{N_P~��|4��_�k�����~�Bm� �d�l�U�r&�V0������$�Kj{��Jj`��@�!����%E��+`��OT��0��ˏ'veQ?xbw�|Y�w���>�kJ���NG��E�� 1�@.[��<�Ѝ76�#<����E�g>�X�]��Oӯz`��i�V�P���+l$����-�u�]޿�r7v
��g��5���՞�2��A�N�����`��yUwڌ|��d.��NF%��G,�����{ y�O-3��g��&��,([�z���^�綅AnSQq�d�z=w���9��G��� 0I�(�94�O�:�a�G*��E�a=��=��"�P��<���� ��X�f��h�f�t�1e���p��a��$k����b��(��r�:�ri%|cG�	�Q�9�� t���XT��JY���N��+�
S^�
�D�l��c�E�HJ �p}�9�g�Q/�wgY�'�D=����2�G�Vz���{�B�r�u�#:���
:sr���ا��1E�L�B�mT�-�`��G@ԓa�
���-�]J�{>��p�F�(N�Hۊ�TC�0��3��,��{����/�8�@�?���NϡD}��O�E-��S��m��7�dP�\"��y���C�)o���=�%��&3�M�*��O�?����]���ZswS��]��'��YH�ֹ/ѱlY�
"�=g���K�e�G7�^�9�1��U��<sr$1�2�I]�� ��&X,x�tն���?�͵�p��]�AřT<C�ʺ�|��8��ʲ�PKCNJ.7L[��:�,[�<�6"���:X����4����'�n_�z���IP0�p����oz������3�mT��8Ǐ���m���n�-r���:��LsGG^���JN�FQS�''{��u�u�XX��6�~��As��\�qL,/P{���z��Ŝ}���.��h_J��/�� |�\-��YM���|T��z���~	��PV��|�� +��s.��䡄��R._�@h�Mgf���2e{���
������hXs��/�i���l�D�L��m�� 0�VA��ޥR"%��h��}s%D�;֦��3\'ӗa�|2jPm�Si�M��ל�����7:��)J��BE�C��b[m��Jpd�����?h����"��,��L�p�p�T3��_�������;�y����i|�w�ʚ{4j�]J�RBQ��\ڥW��^k�r`Up�Oj�����;՝g4
I'hF����xq=�#q3�8�Js�[幁�L�vc��,����ʻ��ՖN�Q�U3J���	�A���I�0ρ�v �������Ӵ�[Nh��E�m�p�A�hON������sh�:�g!�Ep{�]�5!�;j\�^3$n�@�a��>��{{a��f��N0:p0zM�*�AtU�Y!�%�a�����a0�Z"���x=�Ķ���#���&�����\d(?�R�A��E1΄ q��$��'6�66;^r�Pت��Y?�DT�[���S	r������퟈H��1E�޳p�$� ASMӘ<x�T���9c�s+�tg��<��+�ɴLmR��>Н�?������{˕�5��L�������+c��fx25J����z@���b��.��8����	�*���۵����$��T_�/��ݘ�S�7�.{c�n�6�ge�X���7;�hUN���Pm�k�f�\�J�l*���E ��
I�[���n��IM�ّ]f&ja���L��#���{�G���+�A�Ҥ�=^mR;���{����U<bn$��	I'8V�|��<E�5
�/_2�_Xȫ��3�O��ܿ*�¤:Q3̢���~�$~Z)�o�0�w�a �d�ս8��@���4=D���6]Q����/�_�Ԇ���=Cv5~�S�;Q>�#���`����)�|�|Q��:��N�b�
}�,(��o���[�r���iQ��s��7t�$�p�&N[��|g�4��m_Tҫ�Um�>1N����,��&}6p.M8�h��i쵒1�Y����+<��j=t.a�k�k�!H{�g���l��{2�.��L���
:4S�����O�J��iW��IS����V������`�(M������V?�'���*2mE��_#+ڬ�]�����8]Q�}����#�����G�EC��F��N�Q��* ��[q\��p���a�UA����>�P� V�f��N�F���?*�hq������텀��R�-��GDd�>5]��M?P�?J�mZ
��
Z�O��;��rbf�3P�_�E���If1�rd��;��)]@I3�ց� O�m@g�����o+��ٽY_J��6���m�8��.4M���0V��t���@��HV:7���^ai��n�݂�����B�f��]-Te������09��*����_�.�T]#�ޠ�� �O��~j�'�k�����;f�iA8(>j��,���	�6y�Ӱ�T-ݓ�{��_Ǳ$R/ȕ���2�*���-���"X`[������1ɾ���6��c���h�m+��~|O��U���@IB���++�a"҉�ys��HP��?��7@���
�3�4G�8�xB�Q��.�.o)��T��*����|N��P����
1�u~ay IYy
*��X+�ư�ٓ�W='GO�קi���LY�;�Z'\�ׇ��H�+�y2Ro��P��O��ڑ8�l���w�C_�}��a���ޟ)�7�N9m߮�h�!�_cظ�����d�5��&G>7��k{5�u�����MQ�'ᨆ�^.��;�l5;�٢P���0�`gd��d�k���b�H�1�@Ĳ=t|��7=5�j].����k�:p0a,k?����Ԧ��V_98���՟�b���aw9�����Z�B�-pD��5V%ײB�k��2����@P'=�9�/-SG����`�)Jͯ9�,���/pX�����3_��#DH1�8af%q�]9txr�Y�i��Ӝ��d>ř�Q7��_G������%fD0���=s�4�?�)*�Vu�~���w-, D�q?�� ��ڳn̆tf ���+F6�Ӯ�*�4�W[E�t�x0S��m1�l1Xm�&H����	N�2�󮬫�g�j*0�x'(����2��	�p�X"0�(�{0�B���`��&Y���y����08k�[dB��t�)NX�3+��x!L�+ĝC�ǭ�N�͆v��X(�7�tL�+��^[�o�����-�z�U8$�kU	�Ў��?ᨙ�p�ʫ�(�
qi[
dk퓂N >�A�����+�<�g���* ��!�Ʌ8m�F�+��|t�m�Qs�W趥$�t���V:��#�nA��% �aH4�D�o��+U��Rb�ݸI�HU�Ϝ�B�ɓ���ׂ�Y�ǣ�a7��/�[��x1�ֳ�<����3��0�!ڙK=�ݩ�`wG|�! �[�����y�3b����]�JW�OMʐH�������XI� �!�N��EN8��so��(�A����N���1{�J�8�X��_���_ת!V�orUKU�B��g�d�#��dπE�
��u�)��F�W���kث7�D���ŧY��h͢���ʄ�y,���/�j�����ښ��&��C��Lx8 �H��N�St��pi��y)�?wl���
�G�����./�W��d_�g_ )�
g*ӡA�at�b�4јMD�?�%G�*�?�l�}^6��^����^1�E�2JǦ}M2��t��q�.M���Ԁ" �R[�Q-Y�=)g�%��j̊-��`�[-o;�irn����4&q�>� ��f�p9�>/������q�pH���Ky)�;(c�o��?&D���H�]�SS��)�V�fYz*�裑�6���×N�1;B�*�0�9!�m�6sq���n�\��h1�z{���5~�mZ��0�l�˳"R/��3
JZG/~�[[�Td|���K���553r�qa�6�R��Ph,�O�r=���)�-��		0�_���W�Y*
�+� T�(�G]Y��C<�ކ�P�r�<�� �a���+b��{F��[!�]�Kӎ���e�
��1t�D�"@��L�<�����/�H����!��A@}}�f�K_�0=3knM��U1��6��my�q���ѱJ`��JW-�v�ZS�2, ��+SV'��8_=���+�]UY�~��׌f~�eR'�-E���To=bOz��X���gWY���P����g�`D��U�T۩�z ��,�$��0��-�r(*�8 |ܤ��#�vy�R��a�u�v��|N�G�m�T��Εuq��A$@!_��~�b����F $"� L����2�>Sdy9)A��B]�11|X�N�׹>3۴��3���ݍ��vF����{Z�4�A6|���d�vx}��-w����HS�:�fG�rJG���'˿~\4��Y-]e�>���q-b`��8M�{�NA�<�����i��!����&o'�Z�L���)�V���zE�W|�� �` ���BP¬������<��lix���z@�_��e>W5�PA��-���.;�tpS= ��+?өq5�U��+�2���\���k��@wp%0�ۦT}��SL�L�]+R�A��om���L�ڵ�I�h*�A�_i��X7U�
�Lb�!�Z�:/F������� ׳D�9�����4��7�;�&^��%�)���|D}���2-�~���A���dd�ob~�>���)�2�^� �U��j���"�#�T���NE����kK��Q����r!a�N�<��v<-��d���l�C�sᚃz���M�� :�C7��E�Yd|[UZ&&m���\]����u����b��cGdC��j-r=�R�^G%mj�
���7�%��q���6��m��o�Y#�����x�k�:+F�(��~����sc*
\�? ��Au{���9/^�ݔ�V,�8�Î�6.�>�}�����3դE!����m
��]ućE��q��S�����_�U� �R
�h���r-�=�̛h���\~k�W��M�H,<-u�����M��<�,�]������)��{�Q2�S�Mt�Ӆ�PQ�����6���`~!��jl�ﾮi�Ft�m����j?��mͷ�k�$��I@��漊��:���+���ᥰ �T}����r�gM0^��pS�_c���ݤ������-�A��$HIN��	�p+#g �gy"���t��u�#���'����������wZ�