XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4W���o$�Ky��PZ�[���m��ٸ��3+[[/M/�R��=�E5�%�`vP�`�L�XŞ�Ԣ*K����Y��:��ҎG��&�� ���'��4��+
��8��o�bg���C�%׬\����e�A�s���f��m�P���(l=( �Ƙ�6SK�6�}�H�'�d�W�P;%��t٫�1���J��i�xV�\�v���m"��	d>��e,�J��0:�t�A���wB@j��_d�@$g�ŭj���`�|��傔AC%�<TG��H94���"���5ϓU����!�>�j�;���s=��=#i�u\wکA�����)�yM�����37��〸�R�?�$\��Y�T�,�.AR4u�u������6��w���)�^�IIq�y8�*�L/�0�T�?/:�+O��i��ؘ�w�8#qej�r�5%Ð/����/2#>�V�X����Yɘ�����9N2�z�.u��fgxuH��e�L&�~�}��6з8غdv*"\ϝFrC��Mÿ�f�i�F�S�L����R������toog�0���_�SOf �W%>���1��2�LB��>2�M�TV�Le���]�#��O����66,�!��s>
�r�u����YQ%������c�o|�5�Xx*>m��9��"GZM��;��_ю�ʾl��u�P���d�(>IN����Q�[��?0�xM��ʹ�Z�.�o�#yj�YGҮMþn��1�&z�!bp��3��XlxVHYEB    fa00    2910������u:�b� �%:)�&�Q�
#�ۧ8�����ӆ���g��ClD~`D�
E=�8\�A�}�1���E���вF���Q>�H�5J*%n������>�d᪒�Bܛ(������D*̸���2t݋;�]M�|8���̩�1�!�h]u����g&��zT	�����)Iy`��ck8��9��E��f�s<!�����g�翕
�8*���H� Z��Ȏ��C]]�XiY��D�^���6X�Yye�5ǳ�5d�p�r��[�G��7�&��D�F��1~�����0��-�n;@j�p���dU��RGUś�w|
]�5'h
�,f�=ـ�n�%0�����}+��#z���w��-�Ol�L�j�m
��̫H�,���uG�^�\�dg��4�; ��w`q��ӀY�jવ\�mg0+d�:�k}�2X~�þ~�&SX�׵�����TA�ܖ����k��Z���p2=�H����c�b{�rD *N�\8ؒ�G�j�ť �,K�T�6����$����k8W�m��a�#�kx\�!��c�wӏ�ICuYc螂�_��
{���GÒ*��o����jS"�JT�C���|����c�Q�V��@P!�&�R�N�^Y���H>RQQ�DP��_/�� �e^�ݲt�� �e�_�u��LxNˑ�g�5�Wx�CE��<G���b8������ƀ#[O���S//��Y؍Pz����H��{v/3��b�|��ݖ�<5��n�kgK)�d��+���*ʃ`���0q����J�<�"~�ci"�'BLkY6R���~�⌘x�V9o@2jN%H&������9c;�k�h�MuA)_�D�ܨ�`F?U:���G�`pi���IJ���I�S�7Q������<}�33��dbLc��	�*ϸ�[���f���b�~���#�;���*��Q�}��3}�xk�f���7���P�W��D�Cc̵�� �� W\%󑶴���I8�3���A8$侴�Ȋ{����pj������"�w`�gCc�6k�C[�<;͜�F�b��4ome�j�/4͙ $��C�B)�7و�d�#ۦT������R<ڎ!�j�4¢�@Ʈr�$-f��`c��(�8೐Z��KjI�<��� �0�$|�A��A��5S-.�W+[�s�{�?�)3�|%����h6���*a��vy�Y��p6Z�a�0	w?�y	�tQ�,��ƮO��Е�	�L!l�ڿ~�[a��K�(��|�-�Hd ��v�׉ڌ9c\z���x�G�W2�`{@�1�g�H�~�$�dm���_�o�)�~؁�8��v��=r�B(�n�-�公6��j��_�}?�u-E��A�[&ZkW�vM�{}���+cz�0���iͷ�-iliM�NX�hv�>�+ĠQ�N�h�c�8�CA]j�]����F�|���P��wy�2����<-�0@�Ц%�w^����0M��Y�2�pI$Z3��L������(����+�~2�	�<��ܰCk"i�$�+{��&ޮ"�UEkd�>h7s�r�-�:�<`	�E;΋�uy5R��1���Yጬ6�eG^䦉4�؋�.I�(˞��(yϛ�l�m��J��]�ƹ�jE4(���ګ��/�Q�Zא��.fb�E��_v��_�.7R�T*;��e-�B�&�J}�e:$n�+��K���%�ꏰ1�tW7��JY
z�Ȥ[B�X�f��7M��A-��y4V�W��E7�lj��-~��Q�d<�z��m��E�*��@��qv-ISł[߉��5]{�#_���^�ȝ�nY��\񹭎��*��-��(��._�	8T�6�cs��쏢��z3��o����Y |�Z�IF����6[�VL5�	�Z��^�摕����bYM�0?���} }�gZ[���?�/��Q�Nvq���]k�d�BJ��B�������U�G����A;E-�t��8���	bߵ+��ۮ~z%�\�ʑ��.o�ޢ�����w���j��l�MGJ�	�hU38
�WX�8��0�p�:Ww�"����n9:�qƫ�Y{0-��w1��.	��^g.��먟݁������o��4>�V0G �c����$��w`��[v;���
o��麮K �t�(�3f�����������q�p�\l��Ԃc۔������	���t����v�ʯ�m^�b��T�RIao!!;�.�&"+�Y������X�<��W*P�Z��3F���(��O��qw�hāP��]j�9{�L�����%Q��&H�^v�1���xo���垻�کz�u�;��D��!�+|�I5�wny����z����c�$*�C,�_��^��H���KjJ�fO�{�����?����c�"5!ؑ�����(�%'�_��##�He�9��_S�������<��TV<=��h�䒲�,�/YT&v����R��$y%Sv����I�`}��ţ����CL��w@ )�b%jB�Jo����6��E�R8B޷3�'
�k!Z�:����h����NF��p�W�[9��G�	D�z+�M9�Z��v,�ӹ4���Y[P�Uf{;A�� W��k@���%�9Ǭ],�8�j�Hfґ� �w"tљ{3���#5�`�]�GSw���V��ٿm�čO=Ԡ>OF�1W=�X+���-C�qN�d��ԕ��N{WeM���?ƤyK-����ć�4����{`|�DQ��d�(g`�{�+��ƥ�x���n����P��hy�#�w����.x��W�0:��G�|�h�@����|�K�j r��?�k�O���o?�ɫ��"~(Tʒ
t>/)qN��&���0��X�j�4*��������3��I��,5�\R�HV�tE�t�+�A����DIh��GX~`lT ����,�%�8޶ha<�c�,�kpP&ܴ�l�La�,7e��U�l���y�A%5Bc�8��� PĳF�SLszX["��L>/	�a'����\C��!� a ���Y�A�24Ԯ^Dk�y�H������5�� �%�:F��S��#p�Z�ո���ݘ~Ci�+ay��^�H.w!u�\�^PdS�(T懣Ĕ{5��'��vqAn��*�ϐ:�}����!�2�H�,��e"~��*�G4��X�J����K�ĭ�<�������� s�9/k6m�N>6�������|���(��}�~gH��CI`�'���ʷV��A�D�x~(�`jFj�P�1E|�2bC2i��6o@�֍��q�abu���m��/,��8f��x�Qb'������(���N��)�*�cXj�VgS������`n��J1�c�����6�7gp��$�?��a��l��+�䂼k���&����c�=�S5�K��[�)=R�/j�u/�# 0x��
���<����@zwq3���v��{�=�p��8�T�hP|l�A��qZɍLb��3�!Y��Q��,�r�neT��"4�O�&p���pW�v�N\�o�D.�"Q��d��س�-F C�⣥�Z�࿑d��zi,C���Zg�|K�tٍir}~��qzpD��f�(�9qud��e'��Q]d�/��i �R�_�&�V��;���c�S�Ѐ� �����Ӓ���?�qJ��v@;��-�	.��c{�i8!rI*��i��Q	��9��Θ�P6j�Z����_�2-�m!������l)Lc�[��|��\�ϒa"o B�dݎ�n�y5�y�j燽����C���5�˔u��(a.k|X��K���8(i4���-��!�N�W��~!�����K��,q�@�[ ,9%�(�����x��p�Kp���n���l��H<ox5��gj�c��?�v�fa8fy�q�5���?�/+�RS�"��'z�j�J��?���Kg��m�C�=?���ڠWG��q�݆���J�q��J�]Ok��TaM���!� $�>h�3b���R����h���F��c�k��EŚ�g&gmA.���~`�{8:��4��2O<{);2*��w�:v����j���O���GЗB�(X\��*
���p��@]�����(R'��ߧE+n��|��]�M'�����ЍF���`���[X4��41jvȗ��oLH0^=����E�"Lj� z0���T|�򨤙�1�;h��E��n����B�ād��x5,��ˮ�V�j�#z��_��C]J(������PoA����n��#�wn10���j4f����M�S�	�-�����)��f-�����>�VC�W��t�˫]Bk��*%����h� U�.�oÉ��P�8E�ϯ��&��˾��)��'C$	����b������3v���(��O�ꇥ��1��D���(@�v�{�T����R��e�L���}���-�r�`)�5�������B���2-�N��R�*l��oBʷ@FIhC�2���`q�O�]��a	]�fH�f��VR�m�_�k�9�V�(` R�/�h�ƻ Bt��W��Q��^C'����\tIj��!ң�Ͽf���u�u��?�K��Sj���IL��{�-g�DM��'b��	6ءx��0���׀����"�[�&��V�%$~�"�/��'��'��QxӚ�	:V}�{��T���C̰����ۛ�����K_VSJus�g[	_���a-f�#����4YG�F,��@W�\ҁ!�᳀��)�q��g��n�d��+p�R��p��Sg��٫��5oar$��xs�yFMbR�+a/g�R�I��Uބ�a�B1�u�4�[����E���>�GX~��$�E.�C��97�#��,E���pY��m]m�n�~�\�)����+�ȅ��2�vŵ�N��#�iD���}��3d�@4���~��*�*�"P;���@�H,6��uw�������+jNQ��g���_�n��c�bs�T�;T�{l��]z?�(� с��ۡ�_�n�&Jh|c�T��@���G�!/�T�N�5�:�&)�>�u��ꖪ6��x�z]s�u����pjR�����mX�{f<je�SBJ߁Q�s�7����ܧ������Յ�`u�� �$V?1g=�����q7Vu�C���*tϋ~����̻�fצ'�?&�����LYWJ���iD����Gs��Q,�,?Xg�Y���Z��Bݡ�=�0̟��@h2���NY>Pj�,œ�Ko�L(��/q�M����}��3�Vj'8��z���j�P�*�W�U��L<"�.8�T:�ry�&�Yc�gD���>%�8Ƃ�ey��u�ޱ!�'ʡA�����%.�/�[��g�TϢ�dcOۦ�jm���y;�`�#��k�|&*a������dH׻n"rj�VV0�5��e�*��ؕ�A���wI2��b�J�kME	Az��(jb�B�����z��= �ޏ�s[$�	��-g�$�p�}����2��.���f��o���'3c%�D`��K��Ǡ.Jn�^X	��QJ�F�D)N`���>�,��3	u�s���R=��Cj(m �Y�/�nk
+���k1e~���.�.�畐��(a�\�bk_�@�=^��A��舾\A��g�Q��4gT��UK�e6d.�����ya֍m2o5e�(9���28��J��q��%���Q֖��y����xM=)T��5av�v�ym;����� �����q��&P�]�ʪ�\�'�g��"� �%��#�8�߰:�5�2&����]�h|t\���u�������(�ظ�M]�46�oT�1Xf��TzRK�
V��������\��r����j�xǇ�m!�d���[��Y�I ^��v��;�l�1Se9���vv���ZF�?ð[�h��Ќ�GD����2�Uc��Ĥ|��6SZ3Q�<!�סּ����h�w N��8`�ו1�?���`>;sn?���ā[���K�8ִ�V�4�:y�uވ��L�7r/�K��^��_$��9����7�8��"�]�C���/*y���40ȥ&ӕ+F�P�)��h�D&ϩ5�<�)T}~g[w\����h�맭
L���%�p�q=���:�Kv4���{��z���B����L{��òw�\kf4��2�<��
����f�~�ʧY(���r>�b����ɸX�q�f�㱩�nK��b�rL8{�/,��^��n��HL�>���s%	l�j�5��fh�K����T	f����tI�t����q�P/:�	�`�s��+���4*�v�p�q#o^^ӷ����	0�X�A,Ň-�y������V��d!��f*�Dp���@r~��C�
�y5X�O���>LT����[��5���Y.�^���t�[㤎��z��������-�܈zȥ��W�VS�z�������)6���s���K�yI@��{�w��omjo�q nS�!�57����M:����/ے�{}�G{2�\N���X��,
��k��\5��F�P�d�A����r�%�(��.]I;���]ҋ� ����Y���L�`۠�n��ۦ8�v��Ep�>C��[�����w�F�;n:<xH�(�[C��:���Xp�D�[�U�ƶ�g�Nٵ��Mm/��yk���y�H!���#7��D�O��?	QQ�6s�{�M�ql����K�zC��Xͭ�n!Z�����N���)��aB[Ԅ�I9���֠�k�_��4�L^(C���OA�F^[��E�(���,b��Ƭ���>@���9K�)��!���>�˾��,��ٛ���S�H�g����=�6����O�KgC��g��_܆��F����h�(!��f���^�Q�&��h$c�`��ks�^����-ֲ-�����[�=e�cY�=��M�	�!~i Ei3)o-�f�p����BU縩�#�|Y\�x��Zr�⏺?��xGd��ߤK�ɫ)� ��|��Li�$քW��Re�5R��L|���U!+�-<Da�y&�H,�l�6��q}��s�M�_��{)�V^�HR��%JS�J�̃�^i��}B�/6���z ���@,I��@ٌ���k���i/^M|�<QǓ�!r������K`]Vh�*��̼���e4��jD�3�V�A�#�*�8utO%��ﱎ�}(ـ�#�� ;&=T�~�?�:	z��{�
Z��󰏲�;фD��k���BRUw���R�Y]TI����:��9�\FW�z�*'�I�U���&"�;up0�3�`�+},���"��k���ѹl�i�)���U���x�����м�ƹ�d,�0���v��A){�<�^,���g��}[sj^��/�Yt��[LHpw�T�#��:`ݤ���%��\X4T�1=�2sF��2@�̴%�ω�D���'#v�g���-���Z�^�S׉{��ܩM5(�V�O�]��PW�4�9y�G���Q[.���u��f�f:�/$���5��Nׁ����Db�����ٛj�Q ���$T�r+B�&v�8L�FD�ط�A���=�I;&nM�Y�`hz�#�}ޥƫ��e[��ܗ>vo!�8�$.>�#A}"��zwc�<q�j/Ai�='��K����,.��|�l�����m��̄��W��i=� �Vh��w�:����{Y�+�����Ƀ�"-K�/�߬{�j!��E�s�x?�78��Ĭ����Z)r���Ģ�3�B�5����}��m���������1�ݹ݀�,������s�����{.W}ک����m�I�jdm`d��\��<~|��LUr}"�_f^R{���ל7�ޓ!����	92�'�_Kl�OH�k�a��l����o��,��w�>���L�m���>cRU��ta�"�Ã��ڜ���N�e��O�|�Z���Fv���-��	'�FrB�rQ����G�!a�d��r�Λò�|:����1�Nl�dS&�?��@�}��2���&�'��	r�-�F�G4�i�*݋��"-�$��v�gJ�G؂ ��V�@Ob"8�~�3c^9�Wi`!�GǒWH�����#�=:���@:w3�L2TQ�_0c��ƾ�ŷ��[I��5*^*E��G���{#6ʚ��d��n�TS�A�m�����&��K%O/�5;�`�[G�5�ܯFl���a��E�!w'�)t��ɔi�&.Ǌ|i�	�Z�I;\�p��@�ۂ�]ݺ�=��Rm r���p	��U�IM�.���TI���۬���G[�� �1�X�.���w?�[rUז%���.��$�fj�(�� ��,Vȿ!�k����z}(p	�|��֮MVHxf����6���޴qDMO���P�1��}������oW�!}�19Uf�v���'��`<<�3��p�����t�VjR���T�^qWY�F�ڋl�/�А��lԍ�;pƶ2;��6,�9!��j:|��@3tA��4�k"n�9a���<�`}@4�ы���LA	^Me�*�$3+�;�u�����n����.���ö �<�mȫ���ڀ$��p�t��1c�$B/X�D�z�=�|Au��EH?*�f�~�e�TM'[��L-f4>��׿�`>�s���>�����������!��[�&?��.�B3����#�)���ZztH&��A�H�`<a+ZY�[�ɗ��у�Lpjd7�S4���_�'� hDJYܓI���ng+���:�%mv	}�K?���i�n�����)fս��7�[���yj��.�*�F2m�Gp�Ta~����vA�u�2�p�Ǒ\%m!��GwĖO�U}���h�n��
��J��&���P�i�>e�#d��4�le2�`[[ќ#!��:2;��\�����h�Q;ܷM����"p&�`�0��4��A�*���V��y��-�(�X
�����t�Pl~�Kj̀�TԂ��N���y[�?%����뿠{ܶ��E��Ls80�H�7ב�
��̻(�.�oЬb�v �����za�I<�st���A5[��OQ �i����W�g�Yxe�T)�(�:mm�8�'���J:��F��7SϤ�w)�r8.<�h� �����&����ޥ��e��Oee9�p[�;E���.�͎Ĩ����T���c��<���m{�*!�8��H>�p0.Wl��y�t��Uc�?|ӲLg���|0G��zi� �p����C��(�Z��q������[��&���B�.j�|ع���f���,�g�Gi\����ZH;
ucx��������ýBŴ�/��<�i�Ϸ�lo����Z(j�0IPn#�vZH?��&�Tk5���i�^��7�I�c���.�^�q�;!>���{�ks:�1���o<L�:��و��u�u�D��~�/+u��s��-���
N��=E�,�g��&���Q� �Y����Sț���'��Ĳ��4[�ą��Z�����$��k�dä~N�z�i�F'�
���ўl&ѩ�W8�M{�j^�u g����A��*��H�/�����Փ�b\�g������@���J:�{���غoA�{&moN�t�CaԜ A�~���;��qu.�Q!9���quC��l��@�d�*Zp�Lv�3��)�9�0D�[��ʿ��b�v�a�5���������+$�����#٬�I���{�m'���s�-N81/Z�
�2�Y��&��o9�E�dInd��^_�������]w3�]��[V-ML)��)#GjIo0����5���πƳ���A�zJIcXH����}j߆q�>�}�*Bq.��W����/}�T1����̻���i%�|��k��븎c����t�1�����ם�'	�����Y���X�rv5jHY���?�A��'���j\n���V��Ub!���'�� ��J'�ƂIP�Laׂ��C�������P�+�~NW9�''�Ⱦ�$e3�����C��ɨI���B �;dI�Q�
tʶJ.[)�Q��,rA�#{"b���q� OP O�Wm����A'�8;�����@��@��YI����a*
ە��HÆJ,$�H����¡��U�i���5�045CUL�.�껡@(�0��d!\��͌��%+���<.�����|֨�����W�~��S��j{�#ǃ�4�!���,clmR��V*�k:��񨏯=��tܓ?���oL��}�2ZT�J�%�?���]d�{��Ӓ���@!nU�=��;�[gљ#`�[? 	3늴�֯r�q�h��n�lx�X?�B��+�\��ڬ�f;��iS>��*D
5�J�<|��hmG��d=)		�ȗ�F�䌏����4#]�O$b��n�ݐ�Ԛ[��옐d�h���j�@��l���[Ň�2g��F bdc�j�C�%�HΪ��.�XlxVHYEB    6184     f80�<�MZ�h��<��5�lCo�+�4B��:��iaZ*�x\Պ�孈��ؘ�.��<X[[��N>��l"��C9������AAAN�B<	��
��'_����|����^w���Y�Fb`e�n��JY��Oy5��L��]��l��/���И�Z;^4[� �^8nM��/��G�#6�h�،ulA �P��h����>�Ĉ�{�1/��&�R_g��l�Lg�d5��܄,�x��f=���a�dN7bp:�r�Z+��b�NIiM
���`��b"�v]�[�v����.u�A3ޢ�o1��}\�;�&�Ӳ�}ң��dS �ר~ʵ��r�yI�`�zMJ\_L,=��v�7<ߡ E���I
7���b��$a{���h#^���%���O�n��i>!� "h��e}-���:�g�̂&jn���$%߂U�6B|�=b~�v�&|0R�$�
B]Xc8t.
l%l!gp ��z�y0s'%!�Md銽9�{���7Rh?��7o��2�e�"��y�`*�]b)�%�#����b���3u�=Ԃ�ѐ(�(`�F|x'���'��AN L����=�dl��&��=Ee��IcUny��� �M#�~�J&��XF��V=� |�f8Sc=ř���h9�� ̟b����*jq./j�r���O�ZK��.�Z�I�̬5�4K�P}�����8YDI�xτN�)��Ǆ�}_�1���~�K�,cI6H:0J�lO�>����NNwI�p4	�3f�� ��~�$�9Z�0+���%'<mZԳ�i�� :��=���
�������:0�jۻ����R�<��y��X�+���a���|�4@`����ܐ�=�nߪ��E7/���S?p:$c��4>�N��<�\;��%�R۝��wӓ��U��ߙk���S�c�(�"
�y�� �Y
�z�t��x�i�Pb�}�$��겦�/s�r,Y��)tdq�G��s,S��/��Jˏs���($"�����p�9�|�Y�CcԸ��7$����Ni����c����Q&|�M����Ƀ/��K��M�v2�
tE(���jN˰������1O�Z�Y�G|\�����b���C�(��E�T��/=�C*�G�k�!~;��Msg9�_?+D�A/+r��WnY�#�_�3"4!F.�(gPi�w��l���QzE��S����@��Vu���ʺ@"�Ney�Y�O�#��Ɉ�oB���dlqH��s�uz��Rµ>��a 0�59m��շ65׾��6�R��6(���m(Kw�=���Gl��%\Lug��tJ�A��D��0��6������Y�_1���Ík�uBSw6�T�3��\}�����T�=`�O�W��c��Ѐ�?�7<rk���ϭ�o&��a���}���*�0���Z���$����JΨ��`�v.���\Z����)������f�h_Cd�k�p/��D���RY	$��6��hOf�G
s����-�����>�6ؽ�M��'q>9(�i�5S��,S�}\	��X6�Y��H����f1�96!��wL��#�rI�}W�ε��i����~i���k�2�#�e��z@��̈`od�S뼀 $�z��A�#Ѿ�l$��t%������(������)�W��;X���"d�{���j�o��`�X{��˚�9��|s�2�&l@P�2����ɔRk�5e�8�(8����e=��P(;�
[m��E�y�/1iȚ��	0����r*p��C�:�Y�l��r��=��F׻�(��D���BΨ�!�pA��Q���ll�ڤ�Y�P$.��:�?%��ί�� ֻS�(�^-��&�}�U�~�_��BeT����LL���֓�k*@�wz2�:��|��r�i&�H����n��6�p� �ZjBa��D_2WPa��	κ�n�g��'S����	qE�1�By
#_�U	���YD�С�8�QO`�H{��F�������d�f�8���;�[���ywކ�x�:9H�np��?�A#�V�Rҍ�ЎΓg^��17@��c������sG��`�dX9�_�r�g�곍��ڦ�[8峃Z�<Ƹ쓸+�����B�6 <:���+h�n�Є"�.��u�Y���*)����+�?$��;bJ��(&�Q+V�_\�����t�m:i�O!%��Q���Kb΍�~�P���sv�T��*��!^1�g�ˤ�t�IL�DsP� ��
�W^w�`
�������v;(lHdC�/(=*�!��Q�I��k�*��C���/�hu&�(�j��Ic��x��������i�i��� �<�N�YJe�3���5�W�>��Ab<4��q��v�H-p�&�BN���p�~�7�C�,d)��|l���ьC2!51ŏ&^IlRs��hp,�ʅ��5obj�6|V+�Fwc$ �UqH�@�DL�i[g�|����b!~CL:����;f�à~#?P��8���Rr�TԊ�������~����9z��L�l��#OH�)^�׎+����5�?>4M0�8:S��ʗ'xۦ
�?9-�N5{NI����TD�Y���@E��1��G�����bkg���lj$�~�^�k(S@��zm���\W��Cլ���W����"�RC�t=X����BaU�3B]���L~h^�Kɦ���y��'�5l�h;i*�NJz����wj��N�qX�Cq�1]n�6�U\�53����+C�{��e�f��o7���`�J�RF�˔�beSֻ�mO�b�[0��\��@%��_��4B<BLm���eTE.d��e:�o��FXg����٨� ��%\�?��[�%�M�!M����QK���B�.���B�%���X�K]�}+O��{�f��Ô��ݗ���l��:��^��-��P�<
���HE� ]�;Xw��_��Ď�z"��h�Jz�Uic�:`V��J�W�����aў�y܃t�3lmخ���d�?���ű��f׆�p
mok�2/�gN��4uy/�fJ£�UYj�P�O'�,�?�܇���T�|�h�t�">@:��S1������E�'Bwk�B^+�G�B5ۡ�~�B�l"J��N�ly��ݝ�{�`\�(��L/Ms84۾��>o��>���Ť�q��+h0�c��Z�\���ڊ�� e�y�L��ti=�T]�
=�pm??-�����9�!�:���xO�C��Y'����#�Y«���VrA,�TD�/�كԮU>�;�C�`:�]m�;�"WBt��5-�Q�>/I��5���7���xT�	��ʚF��Yb畼[/��"�{�
W����!l;�t	~dl�9��_�U��_zz�4GT}؋�c���S֓�/��-B���t�<��� ����K����"<�M���Kc�WD�9���i����X�+S:�J��D�k�G+�]�h�s��j�ϱ����N��ΩM�
�3*�U�i�G	I�K�P׌�x+���0v�4�~�=+�"/T�]/ 8���T8YL�����X�D������Κ"�i���ʀ6p@+)隺�r1b����me!q��@V�AS��<�;1|��'ێd�'��J5&�^Q� �ƒ��V�W�ęwI<[�����,����uq���A��_���$(���u���>A���+=\e1Om��$<�e���^����^gwkݣ.Upjځ���o�&����^�"�e-�@"�Mb64W�kI#� �T�+�Ġ��%�Y@d�I��;�Ծ����)\x���`��p��b�'w�G}��w�� x���\J����A�AhL2{�<5mf�����-�í2k��	"lbxbỲpa���eU�����M�~�h儂"�4�N�я��ֺ�I��ҀB�BD�G%��2�:fV���	��"�l��os��=V�v�+�o�#����xm�L���|��A