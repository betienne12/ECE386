XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������#`��Y*΄'�����9���{�_��B^������!��V|��nArf��n�䛣R�L��Cw�ǮwKJd����E�#�u��t�����>�~�m�7�YFp�b�x�z���^v0��U罤m�W�K� �p4f:�%�t-
9Ani��ڞ t�=":m���%�\l��4�4tϷ��c�>��Z��Ye=����W�,��O��@q�J�L"����Z6�}h�U��w�M���A�+����V�zQS���Mu���WLI [<3}���\
r��J:>Œoq`w�LmSI,�������tv��c�)���0U�υ	0�$��۽O�o��~+c
W�I�ݘe�!-7bI��o��Zz:�ƍYhu�׸��Y��n�T�����g@Dm�Q��pG���'�iKBچ�=�v�>:	H!lȹ�!�3>�`��R'����,hcZOƅIL��,�/��5�����#$W�J��`�h���R�d;m�zU�91��g>�����J�*��a�8��1`�7�H���+ƚ)mi�Ԑ���Y~�g�]@)7jʈ˒��Ǭ'�z��o�J�7_DVhr�*j{����X�ඈ��ѿ@.2�$IE�T�>�O�a��fa]&�̩���HJ[SO-v�fȩ�s�������@��F��3Ɖ���H�	D;$�!Â��D��U�}CE�b�Zϗ��h���@�L� �n���3���dr1���r���R�?��d
�;�O�P�{4 �L�������CXlxVHYEB    fa00    1950��9�2��F�yv(�%C(}�`yѷv�rڨ����v�w�	�G���	a��]���}�D1�)�C�K�x?s�X� /��K*#Ёn5B����?��41c85���!êWr�~�
�_���5q�i(@����p�<�;�M���ƺ���<��
f�E�����5�g`~�Vm��T!�!����)�U�V{&~w�-{��U���K�{�����u�� T�!ݕެ�P{.U�"ro�7���L#��Y���/1�9t��4�-)0d��8b�av?
$�v\^�,=�1Z����B�h!˩k�w�4�MCۢ=�d�Y��y�t/{��Y��È�]�k��֥�p���M�O��\6^1��D�х�����dzQ�KdjHy�]�N�!Ց[|��߁������nF�K�� "�kù/�yP������p���Q��C~��e�n畬ׇ���G�X��v�㲚�jd�LnY��^��r�Y�GȷEҔ��s4�g��t��+[w����68�����E߷�]�f����@p�53�SV�S�*�eފ�i�w�H�M.U��%���E��L����C!�V��M���!v�p �^0oU�La�j'8�CW`:sV�N1�|�0��<��|�����NѮzޣQ��3������U����=_�-3��B� �>��U��c����xg]�?�6Ra�,ܮQHJ���)
A�Q3�2mw�5��0�hŉ�;<�U���Y>Խ��7�/���.M�ե���Ɛ��2[��H/���mD���S8�$���7��vy���7CWy�V�HI43Ƀz�ϡ�%O�=�Ƨ!�_�Ɠ
�b�0@���Q@�������<?���0/�Ǝ��v"�cy8��@�c����;-V�L;81&��L��X�=��=iQ��#�d�Y���=�=�ꀯ��Ҧ�y���(h�����?��h_��t!���KW�GJ����4������^'��&S�������1ܾ6�\��Q,�}e�4��lv�*g�������]2�\W�i34��*fNJOB??�8B4Lc��uY�7)�6Ń䕣�[=��$V�c;(da�s��+.�7O2�)�`��H��:���1B$YQ���W��
'�����K�\��,��}\��i���)���<Ņ~����Uz�њ����/������"h�YܪQ���'m���0�{�o�f�n'��iYJ|�.���F�V�8���$0���(N` �e�3ؑ�:�}�#�fS���1����¹�J�=`����8�2&R�皸x	�IW�׌�s�~�������yM8J�l$ �����/���%Z��@S�1�_���B�Ex��T��&z�N�З>䳪�h1�D7=�z��Y�^�3�@�h.+��J��4Z� ��xQL$�M�%��٘���;n&�F���0D���3*6E�L��b0W���Z�k��<�u3���n�����t��e<�_6E�a��"#:��߆��l4ĥ�V|�b�j��}����,���<
C�ᓕ#S����6񢿏��]��I��6U2�k�>���!��ڻY�C�I~{'W���zc�-&�%F��'?��NM�S.�H#%��.`�
q�ƿ%� 9В��5uc�A1��C������1+<B�/gڽإ�g��S]
ھE��|}2��M̰#���+r':�Fa5Gh�I]k@�N��G�����Ŏ�������|�����%�Ra�wa�/�[`m�5\��pkb�7J%�F��?���u�IYA����|���tϷ���Д�v9�8��Б�\x���E��f��sͅ�29���P�0J�H}�dp�Մ�B(ē�Q�@�����r��NU�eF����y�R�u�g�X4��q���]9$m(	l�~��j����!̦f�w�ʒ �dVDa���N{��q��#ձ!�y�\B��5�G��9'C|j�!��
k�>��,+�j�����f";��qj�������{���ƥ�&{�0:u�O�]
uS�#� zJ��˚� �B)�k�ѩW��h-	m-�;)�꣫����_��i�e��vc�}�|���=8�S	/nu��T�jE���y�f/s�%��X�詶�u�\^E�7���{ ^	����&z�ۻ��yu��x�@2h�\�7]z�mpHn¼P	m��h�=Bࢲ�G���c�H#�7��k�_���X�]v�ч��֮��zw%���:h�m
[�<0��%�F�+%]�'��ҪM��|٩J��"m80+�Ľ~z
�X׎&ۥ��0���ۓAM��b��S\�N�5�ef�Ɯ������k>f�I}��ߏb��Aw.��O��|�C,����R�Gw�Ʃ������W��f��I/����&57��L������U�����~:����!��w�'�A���	w����aK��Hn���5�֏�p������ܿ��a%�]�Җ���k�T�����ȼ�)���N���9�Ϟ�4�	�q3-���2&�_�<��ϼ��(0IF�%}�2�.mޡ��#⚨+4�u�����{Wº] ��5�!�C�cȸx�v��6ެo��v�F!
c��h�l��/�(Nw1�}�
r�A�Ǹ�"$�:M�j�(#��T��X�d�~�Į��{������f5��-k����E%���#Q�~�[`����}&}J<B"��9�t�,
�7��`s�	QC��9�hQ}p����&XRQm섗�o�'M 3`�c"@��>��B��dP���t���Iw�Fql��>�k~�?!t�I���n�̉��Z�Ž�?���>?H�As��j��k��\�+�5��3���a�~4k�j2pY ����S��I�3&A���#3���ɩv�C�~�3S�Gy�d5K��0j"����y/3�ڇ��Y�����'�1�'�]z[��N��5��X4�Xآ��pJ֠��k�%5�K��*,Ts!Zj�0���,���������
��"�H�G1IzUF��r,h8���!m5��?�嬖ٹEr7*1аZ|\������vu��H���ȫ_gC�N�!ϟ�P�
�S+�/�9ĂHSm�T�
1/&|!�$�"�:���n�}�L�d��H��`}��f�ї�E�,�������q -��.�U���Ó�z�0�ȳex@��[g����B4���Ĺ?q���bOM<�Wy3���_�W�.���9>��BDS�"�O��R�5ɷ��e.�Rtw���kt�8���}�e �2�S$G&M�[��e��T~��E�2����7	dW ��2n(�x3\ab6�d�G*���/��#Ǚeh1~S�f����s_��Z��#��A���=Q_�羫!�zB�Sѭ��~ ��\���<��lꋏ��Ki���)�W�XR{�-e��Uj1���ڙQ^�+�yAG�W��W�z �2��Ն�K�RT%MO��{w�8Z��E��^�~��jQly^�gSۉ4��gu�c����W@�X��*�9M��n�i��C��owYG�(Zߓ솠��V�od�M0_�yu$��cA��d��[mN�����L4�86�o4�I�[��Ƽ����m-���	(gy
'��=��^}]���1&�#X�b��*R��1����2��~S-kݏ���7g����ɞ�\Rt��fe���h6�,�["~���<��\�I$[� ~�ms�8��!�yc������q��2{+�U^Yf.)v��s5��Nm��j��I�����'�lތY��"M����n��d���P�5�� ���B;e��nε3�����yF��S��J7;��CP�GbR��HԘs0�C[��9EJ7o��;)43w�,v��~���+ɓ�=�Mms�9|�Y�S�<��a�F�M���k'j�jH���&gh���n�	O�R�_�cfx���xc�o.�ܜ���{�7��oO=��� ��Ů�!>0��N��\�g?8�d
ݭ$�e'vHk�=�o���C��Η!����0�i�Ǡ1"w�����c\&ړh)���SQ��dIXw��L��!�4��׾z�ŵEsso�m	t��
ғp2�6�{qڙ	�Y��!w\�O���#F��!a5{�U�R��ya癏��$�w�����~<Zԛ�%�7��fSP��(Q���[3�17zXp��s�-�"��ӇtQY�A����R��{�UjJ����ξՂ��Ȑ�i��C�/�X��}�Vx������t��сejS\,{�WmC�9���0d�ƾ�]�H5ZN�9BoA� �f�?J����R!�:lk��Q���E���,���f|8iL���1s?��O2��J�����xz�҆_T�)��؆'���?��ϩ�iN�d�n#*�jZ5l�#K��Wv@�q�B0!#��@�s�[L���Z�)q��T!y�g��ںۣ��2�er�8��WLm����t�|���`=�u����!�4�i>����#�����!�V�/+��C'�t(zW�R��/u�-�n�3�Y�-S�uTL���c��xl3p��0��1g/� J'Cn��,�[�%�2��@�sd�T�������Y���e��7�eɂf�.?쮬���Շ&��	�8��G����Q�^O���4�y�V����(�z�O	�u�rlr%��G���w=��:���y�e�# 
�Ĩ�rL��y,�L�E[V��GfY�`�UEK�=�)���5���K<sbKa2��|�� �k-ht,q�:�9x���gd��j�i�:t��]�S$�M�6�� B��lē��b���L��=���N꾙30�(SP�K��u]���dN��������6�k����2̟;
�O
�{A��E�W�� �*Өjꔀ�g��n_����%{����	����
�w;r21���}SV��.�aխKy-�(�{V"�0@s�J�튵���[�h��x��(��q��^���u��߭��R%SL����J�+���'���^6�`�_cAoPuu�)��eb�]E�&;A��ŉ�d1�B��ì�W@\9��a5�j����c:����q:c���1�*u��J&���$3��پ�ɉ	\,Ǹz𒊴�GĉU/�c�c�r���+G�Ɓ�߲Rk�R����	(}����1ϧ�\ݢs��|�����sB	�!�p�
��Z��
�C����|�(�Ӝ�RF�k)�W�tI���ٙ�w�&2ȅLë���R�Y��0������X�4!RqT�AI����?JPD}	+/���Ug�䰄�L�N?5	�L1�zק��c(6�ǣ��J�d��@��yn����y��*ʫ(��K�_�ᩝ����=Ъ��&4��?�G>��"g�zOa\�"�����N�_?_��(������KZ.$l��R*�@{c1��x,�hs�_�.���Z�Uk:;�ʢ�^a�aD�W���g�:�O�nZ��b��sP����C����~���(�$�j��ms5掅�,t2S�b[j��5��z��ػ���H�iu��/O
�ߤ����"�r���帖�Ѯ�xU������V̫-J���D�bkY�; �eO��p4�������gL�YL��) �Lt�h�O�$��]ˮ�D�"&��ψb��Y� ��~��b���a�,U���o�v���D,���i�m7T��5��_3�1���c�hk/��E{��#$	LC�|㚾<�]�Dƽ*�B�*�l;��'A�яDA�X�(.���vR?t�%�j�g�؂h��J�,�YG k�.��	!���2�J�iB��.\B��{s���1����Muhs�O���0L���~��֦��b�����}��j�	��6���+�5`�w����x�ԛ�����REߕ�9�!����X�-<��ՠ�Q���L(��z�$��������_X�M
(YQ�?%��:�L����w^�am]%���4JɉĿ�g����!w�ϡ&Y���G��H��?�>+\z�LB3�SI��c1�9�g�������v����3ɼ�1�%�[� �ap�v^��4�Ư0Ħ"{ۑ�[%���)m��'8�-0��m��G؞z/�&!T�=���r�A ��P�����mu{!���ִT̈́n�q.V�z�����[2-��l����-�87�k��ųn�������F\#B�k�X6Q�>�D����Ip@#,L
���1@�C���EZ2�ju?8����*�0�.މ=^s���b���l?��d�9�9�s�A�m�}��?Rb��Y�9ːI���q2�1NO=�ERV�Ć��4;�"U&+XlxVHYEB    fa00     700X,Z�9��@)y�)��t�r�^:�fq��
X��ct��7�g]
������k����[��BH_�ӎce8���]�q�e�B|�^5��ƻ.āV���Q��ֆ��B���ℇ�i�BP3�h'V}�I16���<�����ψ�����Z��t��yn���[�{SR���hv��eC�J�GY���:�DQ�\�?�|i�>~i$�}vq�+1T��zn�A;�G��d��'�����Wk,"��V/,�v��y't�U��W��[r=��	9��@g��u#�e���?hn6����C�b���l���f����Eu���`2�Lɠ���{�#�����K��x�מ[e>�v�I�:���8�|x�#]}�~��H Q%I�!���z ��-خ���=�W����dbR"��b2o4(B�w�`�ګ�g)�#����a�ý��8��Ҥ�D��[�Mtb���B�vT��yb�P ��vCI;]��P�6��_�Ƚ��HjO�d��X�7�Pˑ�v`IԱޛ�.f��mt2����>U�yц�;֎/3.n\��$,��Aa|�zu��,�X�`�e���kB��[��zC�DO㞷6�+��h��n�eU4Rd�W�g��_�B���H�k��:.��,�r���ҷ��B����[;��C�b�'w�wP�s�Z\��~d~_vd���*0��m�F�4GQ+��Csu*���T�s�:SA�2�cϯ-'��xN����ݯ�Z5����#g�@s���=�c"6����� ���8�ȨP�	5��IY5��Y���SKUv��]n�&I{11ҷ�ߑ�I��M2�z+Q���i7h�����k��`���4<<6}�ڲ5�ZW���{��eƣY�W��M��v�Y���Y4A����Q��Ud-Ua�jI�C�W�|������+��P��G�g��&�#2W���8I�[���P5����ax;9�����vv��v{A�[�^#E��z΀�¼�^f�ı����~39Z����}���\����.%Ա�7aײI�K
$S(zbi�&~�r/v�='ْ��P�� ;��k�6�+�C�� p�=��&�^��T��!��D0Xq��Z'��zJi�����%ΟB��:�z�;���Z�We1?eӯQII8f0��K�X�[�Z巽�{ϊq���ۼT���&�DfA
]�$=�GY�l�:��)Z~���cIli~j�ǓeM'�0>U�P[>G�f�g'��~;`��z��;�i�[n�#@+���|\Y3���v2!��q靧4��21��y���h.�F5ѧτ��6��$}@k���7 Q9;���^$`wCVpJ AN��Kա�C9p�:f�w��#q�����gCo7F$�͗P��?�6��nBXD���e�%�[m3�a���݇7�ͧD�Л_����y�T8�ᡧGd|���g/H͒�x����~��r������yZ�pZˣQ�@Sy��a�������>0)�����]��ymb[tE:쁶h~A~=Ǹ1���Rq}&Qb�W�㹌�����߯��i��i�����z���I+3� ���{v��0y`�1���8�]4�{�!q�nz���+.X+D	�]/��oO�)�x�uk�7�����䇐~x^�P�╋�<���P�����Q��N",�!��Ѩ�8��)��zy��M�h!I�e焋��`u2�7ѥ�j���@l������_Ӄ�y�>kg��x�J�[� i\�~�S<��h�kEN�GXlxVHYEB    77da     a60��l�6,Ʉ�u�@S��&�V�>KQ�7��������Dl�Є�s��=��P��	��(�|n�z��*qdA�Q�,)��}P�t|�ɔ{�)l=����x7F��8�=!���-[���i��eyD��rj�J��L�V�0����f����J�L�������L@�nR�h��U`�_��25���Ӭ)�5�О� ˾�E`�ϤK��'�
n0��t����ǮW0,���H�\&�@ 2��CC#�5��87����y�O��u6J!9���o��|;؇����_��@�i�[������4� ��`���Qr8k�	Y�+
�J?r�>�E�Evh�PFt�C��g̏�$ '9M!��t��~I~|iAgec��e+�)ם��5� �	�J��$�>��-��������]�R0F�msI{rh+N�PR����)xY��5 U7�П&~��*$4��N� A_��Q^���FĆ>9j�X�����%QϜ �����n%C<HC9pB�?��<?�=���x��2��<�?�ӗ%�6ނ�{����uW�5,[Ǡdxo���g�bPtM����ձ��hJ��&qc��##s��"�{Ģ.�Hg��:fD7�ːk�xX�����P2gD��j�B������|�Ƿ�{�{؈��hs��.ҭ���[���:�K�^�jܑ�.�~��)��(a�o�A\8�XFt�p�[�ڔ��+�w�I5�j[~jX�[i�=�I��|�[-�A����)�� o*��ퟠ|���!#�9��M���������Y���㵿�]�8��u��~5=�	�<*ܧ���!O�L�>�$�2��ڎ���ǰ����S����I�1�D7�%V��W�{#(�>�Qo�,F�tʥD�4h)��Y�̺��ˈ�e`���d���Gc�[�8� fD��a�f�	����.�j�9�>ڰ�*H��+ʿA�>՘F�,7�hK+�p���7�:3_l����!�P^=�^ڑ�`�|�vՁi���t��u�+���Mq��}���t�LK�t(��R+aK���W��|$1[`�)o�7B�}�½m�ѱ�C��2�PD�h	/�����1�t��AI7�T�n� �gG�A>���2���������l]�$����N	�E{��&ɍ"��g�߈���r�(�+�E-ͩ��q���o'�B��'i�؊�~r��Kފ�\�w��??��ʮ��>R�*����P����;���V�����Y�㴚��̽�g�zmz}��\�c��j��ۣͅ5W�OCu1������J�Ȳ˵\�v�?�����0'�r�7,hW]]��϶��"[�ھ�\�u��՚_;�"o�lu�t�qZ�ں���3I|��H����Z���PH��Rc���x[����2h�;��x-�?�eǥ�ZYʴ�hGE���Y~��Б�2�j��/��l�u���;��?�l
i�'�Ea~?�S��9퉆$�����w��(��Hs�˷dm�ag�8�^} ��@�x y{�ڿ��y'����"�2�n᠈s_"X��S�֓L~I�d��w˚F1��*x�y�F��~�ɔ�f�<K�v)p3�׶�� ��:��p`Wہ4�*Ţ�F�񭡣�g�����UQw��F�"+;8�WX��`����)e���������ܤ �5��� <�5V��<�!�ʭ-��TE�O7�I)��P��JR��3�y�4�Xۃi�e+'��K�3Eǃ:��a9�db򱩃�	��d�T��$tQ�f�h{���h
B9@n���S��lU��de���P5J�6ȋ���uqP�����̭��&ſ��?��t���T==�iVw�Do7ͱ λI���l�����b?� ��+�#����>�Jj3�#=�s#�<��P������'_�M��L��%�����Sm+HLs^b̲_ ��|�kr/Gڣ�i���񱕡8Jp�/�� ¼��߂%7��r�=�J:�q覚�E��Dw22]Л���l*Ŭ̱C�`p�� �Ǩ�EَKO�y�Q�N��'�-��p�,��p��̾��F�PX��*P�B�5����X���"Zm�a��Hv9@��XޑfϹR�:��pȶ�O�_$Ym*���>���P��V
���k-��9����Ix��kY*w��#��H�d���Tf�[�X�sU� ӌX�Xi^muW��F\N0��V�~"�)�9ʖ�_�vsu^,�Ⱥe��"���iB��oQ��	�>�Fh�y��_|��YBuit�nq�`:�V
�ҦtW! ��?=q߸h![���s.4m�2�Ƀ��wwu"V�2?�ˈ��F\�J�!���Mw��l��^F [��?{�Y���+�mnF�=�]�r�@��F灐�~�wH�kC��R��'��۷��*}�%��`d����b�Q {��7Q���c�wwW5�@�-�/O�*s�i�Lg����~�)	*�ȉ�+��Ģ裊B���ݜ�³M�����UZ�=��M���2e{4��(4__o��w��N��NQϮ���=�1���|�4�,������X.��s���v`��q�9p	�f�+��n��}����[�{N�����I3ӮJ�KC���L��D	5Ȃ .t&�e�M�ax�