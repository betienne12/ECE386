XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Zˎٟ��2��)xX�*�D
c�<��5�Y�g�iz6�{�*�'7�`�.Enf��/ۀ8x�P�8`������Cn&w�ݬ��[��<��'��fT���G�(��Y�ni�p��[ĩ� 3�	������������l�'H��?� �!Ŵr`I2� V+�*U��^ճ"yf{��38�N!	�0V�Z%ڼ�z!�<���P������2�
x��o
Zcik�\�Og�i�Q�G�3�m_���g�{>�1�ymڶֿ���{�v��yg�7Ʊ����M_�B�YN"�3��Uf�j�ame����͈Β�n~<L�/����u��U1{ދa9���C3�6�]J�V�`�K��vLk�|��Уj��KӖ�H�������)�A����皞'?�d×0���^&j����F��4��ٝL㌻;"�2>�aX�p�\�&�K�GԆ�ۉ�i}�av�j��Kh����B��%����Mް��}�3�����ֈ�Պ
i�)-����k�-��0��97��Tm�5�5Kdȍ�t:�]���	�f��O�5�<��!p�K����meݲu���7�0��E�ր�s�������Cm����<yWC:���
U�霣�#�W�"���L�y7#K�Tr��������G-��2#Bn�8���g���T�hő�$՞(��%���$���P�
�`zPDM*wT�lnԯ..'����"��Jؗ"�����a.�uQ���L頂�Y��*����iXlxVHYEB    3042     c80�2GK��lA���^q�Rom��3h��4��@��K�"����@=��ސ�%�R�:�����t3� r�.�_)�Q)��Ǿ����ܘ~ z�@;�����W�+7yCh��%�v����4��'u����)y|7�G�ę%��C�{l"���>2��I��i*�!�+�I>�| s$�啌�O��}�0IW�D���o�&b�+��Aa�b���WbU���Z�Laݤ\�>�y�Nξ�p�i��%_2�$|�E9;�����54����;�-h�lBi4h���Hv�(���%�,J���dy}����3p��_�>��R=��Y�����!����p阸��0�(��H�Gr��OpP(0�b?/�s�9��jn���T��OD4xxx�J0�_�,�i2_���'��@,��尥YЎ��#:�Bm��Ld;F��&A~3� qI6-�
��"�E���4��H�=w�ߤ�~�B�L7�V�h5Ӓ|��F������⭭~��^U]�؈P�7���3�G˅����C�RKX��sە��BU�ڔ{� �=�?̋�]�`ԭ���`���i�Ͻ�ŕ��vB1{�$�B���ĳ�ͅ1Έ�>w���H%�A�^09�h�N�C<)g:����20���6�ʵK�~%�X)���P%mM�F�MZg/�'$q�u�R7C��J�2s�K��P��5�&G"ƣ��u�����O���E,@&�#�U~���-	n��J�{�\�X�g�)苔��m0�5�dN�":�cy��}�c��mB߲6q����rR��(0YҸ�gG�+xc��P�[���}��M$@�n�ͻ�?�V�B^w���GjA���o���tOEoh)�Yx�^�����H�0�o��ys�4s��Ih�@�$��χ�ܦz�D��BfG���p"�����٬���>��+�>&Ju*U�6	�R����:-+�ULW���5�ݥ�� �⾣a�N3cst��H�m�~lV	wL
��𲑡��a�X
[�9Ǉ��[ou$�t�w�ט��8Y�2bvݛqYzmt�x�#�%Q��#v��fW�M�%;߈�����Ls�C�Gi��c�����f=Y�d]�Wx�L*��>�AˊR��������T�0sa$���.���q�	�M��S��>8k�q��!k�F���x��!U) ͡n�ZX<8R̐�h4KO�ψ3����T��Z��xk=�璍+���v���W�����4��+�)
Y3U{Q/�k"y֋�d���Y�Y��<��:�r"g��>r�B����=�ŞT����.�ɋ͗ �^����>VS6#��DF%��6�Aۜ�8]	��Иh#�9J��:�0CC�lR����j���9�i�K(:��n[d�ŅQ�)�����t��09�~�P�ؔ���v���v��ⱡl��]��=����"2�ϔ�1g��'Q��?���CE�;Bp���'1ʂ��Ȍ�daG[<mCs�a؋>"���ڛǊ����w=�)u������d�s���ϣ�7�}�Ŗަ�0Y�%B'f?`�s�h�U?#t�br�i�owu,5(�n��|S�A��;�iR�ɡ��H0��%B�z**��T�5�g�+ZӹGm���Dl�ls�����	��Ҭ��o{�&::�Q��5My1�����-�y�B�����V��Ց�LdeNı�9Ŀ7	}{�	~!��7/�4���k,�8b���wEkV��I�ó����L���{��_��?<�K�=U ����GΩ'eŹ�'5K�jy)��I�p&~o��2�aofP�<���K���Ws�[����+�s@䜡i��Kpj�O�Y�	S��o�%*z+��/��N��pٙq�ݲ	6�M^7H���_-P���'l�M*n���.Xm�&��^* _R���Y9�>�/����َ� g��6���	���g�c��[���z������dK'`(�8P)�e��Wo��1�L�K�~�����j�A�9�H�����f�����n�]�C�V�� lk�v� U�OZ��55^���G�(���n9����;1��Ŏ y�!����L05�b���o�/|�j(dr����^ĮV2�,��V8'La�v�?��l�w�퉍f~ۚM���!��&�&\�o�!n؞9Q��z�'��@��f�Wu*(����/∗^�D�&���N�aB;�V9멙�on�m4�'�2�/��^:���M0��R4X�+����LK�.�T�p���Od��]LA�����6��������*��`g� �߷�n�zekcD7v���/lW�J��w̓$�vL��_��$TS�V�yn�^Pr`�����X@��=Ѣ�H���6�3�j����o��3�*�Iıl�҉M�M�7�TYX���U��l��r%V29�������6���J�ap�VZ���Fu5�>��h7X0'�����
X�z�Ƭ�Ц����uL�;�Sh����&=C���f�����GÖ���F�Q�����Q*f�t�jA���M����V#�ྲྀ�\���=���-��g�  �-|�v�<"�^IY[g��l8OgC#�_��}���T���N���3���ݦyG���\%��euhPP���C�2s�x�.S��LQ��Ձ�];��F��pH��z�M�Co]���/���d[*�t�\q�t'�����Mi彭���2<�q�$c��p����;K��V_i	h���ݟ�-�9�BV�5�<��N��>}�(������hI��J��ܠ��(;
�����	6��U�����֮�gh�ts~G9xS�:��?7��IX���Z�[�>p��4#�0?W�Z����q�p��� ˝Hێ�0}�7��G,m#o��*^�;�R���$4����������4��J��t'h�C�D�k@	so��U���?!�jP3�FX�I�)�	="VSPR�Fˁg��%m��@C����;sV(�6p�Q�a,h�z��uW�J�cL��F��V�����=��P`�b��Y}�'�
ױ#����ɵrݞR�FjGZl_���8h��mʅ�|��`�\+�xfg���XH�2�(G�}�`L �~pJ~���S�,�bLZ!���_M��v��0���g����	�cP�k�܁Y$��?��h��J
a=���J