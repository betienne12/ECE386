XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����7�۟-p����oCD�@j��J��6�Q�ܣ9X�ÿB��5�GG��C�uR\�><�bl%��.���]�.��0���^�� 8QJ!P$a���~�ʔ	�p<s���{Oq����S��A�B7Fukj�A@����y#q�ע�HL�p�EX�����}Z����=u5A�WM"In��1�u����sD� q5=?�@n���%�0�S�#t�O_�����uQ\��>�vd��
Cce��	T�G+r|'��B�߽���~o�=Р<�������61�?��@A�Js *��3XG�r���"^o#�Kk���&��9I�(y� ԥ�Cg�8���1�:�ԟd��A8���M�b�Ex��4Gl�U-�5`��M���B���� �$l8�?R�C���,|$�\>�r���4%�rڞ�"�r(�S���.��f��E#���_q�j���%>٢����A�{ک��锰����L��W[߈��cڀdMܰl�=��U�2��^n����zO	��t���/�����^)|���Z2@#SMx�~,i�h�b�|bdS{���xE"뿠'Z��^u���904�R�>'ə�<X���˝��5�lд���G���#/������ض%Z(��Ј+���uh�{�L�|���S�"�n�2y�e�ɦ9�/U��I��Ep���
S_Q�}E�b����U��)��7р�n	IW !�&��ьS�Vu*S��\���z,�4Q�oo2�,�yT:p�c�U�Z�v2XlxVHYEB    c3e8    1d20�3/�Oج�sd���k������8~-�VxT�k_�S���/CҠ�z;�5Uj�Ȋ� n(����%ʼ%���Hj��X48�k���M���܀F�v���SC K�~�)%��f[S&bɀ}RC��(}��c]��B0�탄���(�-�GmC�&Ų�tC�L��V\*$#��
 �W(�Σ����*u�h���v�C�o�}��m��r �z`�1�k�m��"ъ�|��������O�'����I(.a{�L�x�u�"OkB����ȫ�_߼[:,�S��!����XN��"yG���B�v��P^��L��y;`4�Ux֡�6Z܁����M!���z����N�.�2s��ٽ�}{�l��+�C���0�+����z�Ƨ�=���9�@���ڼ�N���	i��1>�ZF�:HF����?$F�`�W�\��5B\��Bn�踢�Y�XTgP���h���B0�l#�Q�c'����ԔҤL:�(����YQ��ܗ�nN}�u�=�n6G���o~օ��_4O��3�O������F�x�k��#���"��?��4}{��G�
�k��o�,&"^V?g��^��L�lI�5]��>�7�ʺr�uX�F*�>�7Us�Ocw�)���8�� �s��`��X� �H�	�a�J�q����Y��~N� lw�C3�$s�
_�u��n�Y�鵍�s؅:ǡ4`�t��&VԱ�oz -����'~{V<t�F�{�XQJv�y����N��Y�Ƃ�N`�}a&5+����ӑ>�t�?(���[2�����cy_�.�k�T3{�Q�7Zg�_z;�O�wMg)��;�L� jK���Q�'���>�;^�UEْ'��!��
�@ֿa�3ʓ_m����#޵$��鯬d��v|��)u�&�V�`�a(l)��E8���zЏ�`���GA����ѱK�>F���� .#�Y?�3"�h�yEL�:��3�r�Gza�p�=��^��i�:�� 
>��gl�ռu�?�+�]�m�x�\�7�%(A��l��A�g�������CRخ�ܷ��vh.���:ҹ�ѥ�{ǥ�:��V��G�]HfWD¸�Av6���%�T��C-�;j�>~�ٵ�*�&+���$�
C��hDv����~�u��Qw����,����{����ᑯ*]�q"��,5�_���6�����t���I��׋����7�����Յ�CI��!2��z�R�xo�O�4'���?�˕<m�����H���<u��brI\hxh�A��[�	������z8<��S,:_�Q]RBa:�4�~��k#y�;Y�zņ\�72��m,�]+�$õ��4v6:�t~��r)��y�YNc�����:��y��^]b�e'd���C���Z6�ϊ� ��]��@+�S`f9	}M]�U�IK��,��¡����r;��?E��1� �i��_�s�ΔU�s�؟P5׌S\L��8�&uU2oiƁ�h��}��Dc�`%�q>}�F�w �Pk�L�<�ȁ�t��p?�����[^�Рd/������'���L�^O�����w_��S�yf'򷌌R�`�����������*�!�����3?<��Re�H^���Z���@6�Is���6�%<" X�⑇���ҍ���隆�aZ��oR���e��Mt"�i'��������� g�mG�R��"x@��E��^�nG͕�yG5I����8��i� ��7x��O�9��I�kAѴ�a��-�_�R�`�=�}ğ�j��to����Vsc��ݼOρb��>D�f�Z2�@��{��R����� f��,\>��z���{�> �z?/4��_"�έ������+�m�ou��BzQt����������ms��u�����5ſ�󶦊�t��";���z����K�mڅ������nתڕ��%y "���$L>�>[�'p�9jj5�(�H�K[\c��:e��ޮ���W����H�P[5��\/y}��Ql���DX�aL��9�v5�t�,)_w�'TG���j�?�ɣ�������a���#���&��}��������=�����{	N$�ͨ����.�V���b��Y���c�Yl�:���t��
!`�6^��4ח��^'�0��z���rC�0��*!�9�����U޶��@��?d��y��|���\��_.�1ܗgӥ�@|�F��,%��!Q�� /)V������I7+,k2E9�r�ZB�� ���=��<		�b~��k� ��C@��76��V����o�t�o�����\?��(������P���~��{��Z�Τ�r#2g��Y4���Ce{!�H���=����sB���=�_h�U��$�<�e���8F�5��tỗE��X������`�>��hx��s�z��iDBX���2c�JwCpfKk��i裧�8�9����V��Lm�Zď��DY����t�4wIG����pd��%�s,ƍ��md���p��SL��q�N���Z�:�?uԣ6����	�*w9˹��RF�!�͚�˨F�w	�azH��϶)��)��?�zI��J��9W� �R�r��	���u8S��]���I�����y���������U/}�g�BI�6�z��bjn�\ �Ǭ�4J�N���2>��B�>�'�C�����Ams�uL@PF]��GC��<%�Cݾ���L#o�'�ꪴ�>�x�,��n�Jb
V>p��Q��H�r7xT0��M�nP�h�<�E,�9M�f�e	����L����]5-��>q������`�~B�h�k��?���d�����)�&xd�'w&�l�����wQ/UWD;Jm�$�|��yr�W�n�(HmRL�Z��8i���dX�r#葼�q��N�1��}�]L ��'0��0�Q�p;���C�����k�FȜج�7wD�z�'1��Y�8h�9�qG+��R\�ٞ*���j�;��M�J�����\_c{��?H�P<#��$��� �_7E�=m��g|�ڿ���X��j��rxΒj���l^4�L�J�PHva!�c�B>
8g�(^c]�S��z��Q�z)̹�+B���{DM&�.)֥�@$bO���1"�F����(�˳+2��Y����R�
H� �\#(1N$+���!����`nh>A��F����u${����.t�PO�E�d����Ԓ}�ϩ�0�IQKm��0�~�u�L��c$`���S7�נJě-���3u��UB����Xe)����:��)�Y�䆑�y��^��Pq�5(�=��t�KyB�2�������ˬ��8و�34��R�<i6�('ĕ�Fq
O�/䢘����=k���B��T���]~��ڵ��X�q-=:�������M)\�K��Tm�sD	uj�*,*�Ԉ{"�r�ˆd0ZHJ��5�ܮ8���P(��cB�������A.��W��1pG�|<�t�����2 �jqR��-�&B�� :��1�� �8�o.<[�of�aE$h۪TX2��d��ѻg^�[���<l�T#HY��Pږ���{�댝
������N��ɽ|J"��u��A��NZ'Y3�.
��]��1{��IB���ʽJ��
��̮�>�˱��_I2�C.��J9�6e�,�>��߻@���2������&�V�P5�Ie:���`��9۫�x��fTwy��{�}Ro3�L4��%	\�7�ъF+�D崙���+->�^Tnz�nc�|h��O#	�K%�٫37�0���$4O�,Zv8 a�g����O�n�*�P8Z\�1�ޝN�0��t렶��]>Txw�Y	P��n��# �Ai�ܡ{�3���|Z��6g5�d�a���1�Nz��)�r#|�.mŅ/���3N���<Ow�H���!�r��q�Ƿ7S��7��Tb!���)}���Lc�j��.��P��&����3���<>qt��6X�"Wc�<zj�
ۂ<f`�|6�t��mQ�h(Bh;C�awt�9|�|�}ژ�aaе����WX5>�v�/��71d<�0+�oZ,�7-��1��ɺġ�r�g�g�HWL����%�jc�0��Q���� dfN=j��6nt��#י��#��� x�vR��ܹ�v�WF����)
�ޤr:J�A&	f��t��R,�A��@h2\I�J�`���T i�T�Qn(Pr�y'a�5��q�܊��.y>�@��t�ʎ(��:c.��R�)��������s��]<���SxIK���/��`���4�ю9v�]�BX�k~5R/؁�{��NS�u�(�5��1���i8�hY�(7%�f(��b"��3^9_#��
�-g8�Jk����R���o8�Mؾ�2����<�*�4˛Z}��B����<�N��W�B)#Iw���@Qi�v�E�6����
�wU��mw7ME�'�p\��r�cRA�R�N9��׼��
i�۷ Ѫ6����v��UD�Sɚr�����ٛ�/L�,Ye��O�5��Ѵ�رb-�������n�,8���p���dnXF�k��߈���,L��`�y-WR
��w�"IB���r��1���a���ho�-څXĆ8I����oj�l8��Bu�Yi��J�d�!`��_���`KJ6�n��"KT�
��`({1���5��H����\�'�����D���{"j�[+���P>BT���W����i@�l�6��3�%KF�:jv�4��^����3��Ǯ&^���;�-��d�l���}��̬��@P3Ȉ�ȣ�t�iC�i$	>��#��W��p0�����zD��'@l�vYb�ϗv9�c�ɚ$�&%--z��U!@K��~�M]g�D��:z���>䪕C�}·
����D���6!�-�K��m��O}B��|����!���߭|t��@c�i��������>)�����?�Wg�cs�c�f�B�(.6<t��{�	a`� sZ2c7t�GA����%�����k��}2�'�F2�$��Gk!/=Y���+���p�G�8O�u5���U�t�	kՄl����4Q j�=���#Z��i��>vy���9��E�4���ߵ��)���^`�㵶�0�Jp�DOE�n���C^��/�͏0M�9�NuX�;R�٩�<�B�2n� |��!?�H����0��Gr=�T��������ܰ�h�gT�{j�셃P5Rʬ Jr����R��cҺ���k��D
н�Ӧ��X!E��$�����,+&[X�T�H5=���2��t�>,庨��	c�
�-r��%^L'�/z��`�n%�����4�p�}R�mDEw��-�����R�[>K��+mЋ.2��~�cI!i�_�V�f�X��DA��a��ג��XI�=`�+hW�g 	z����,崴����Z"�z���@Ĉ�es���j�jU���鿓���"�"��YK0G��n�ґ�n����S�z��)��mC�vN��Vv��~g��Z^�Qiv]�u���ū�g*ѯ�}B� �����:d�����_���y�>���{8siíJ�
���tK�`T���N��OW[��v��TXc|��|��K5���R��b����a�4��	X�D<�u���H�7UR]a��~�������Fʂ���8[K5��8���ȤJ-#IY�M��ɐ�\q?᧳	N��W�7k"�(v�0��X�t��	%'���p"�)5kHVx�P�9q���z�!��2yՠ�Q !$@Y����B������ p�^����X?#��G�G�|����~�k`E�<CŻ�HN��w1]6�+�{_&�!7ĘG�Sb�]��BlnV2�2c�JXQ*�@��&Z�qg�׀2;dXi1	�0.@��gH��$׎i�%��м|*�i~3Q��#?�"�3����m(M�V����]̖0���c�rg5�����Je��W+|�%tˀ�𺒀5K)��V��Z�"�}d�W#������ �e���ܬ]ֶ�%����� �?����:���uo����B��ۜ��5k����>ˎ��?�qԁ�Y���*�{Q�+�x��޵>3�(o�X�<������&����L$����������!`��'
JƬ4G5�/|��e���D����y>�p?J����d�&ކ�Hw d��p��h!Dl�\W���w����}����A�0��d�F�6�P�T��=:�U�r���m�#�g�98�ҙ	.�th}H�C�wn%A&�{��.�1$��:�dT���S�@@̽��wlr�� �-�_`$9�Z	�2����Z�@n���;���p����璜��4FѪDY��at�-�d�⓿��{q[��g��0�@3��H���ي(,x��E�2�qꝔcq��IӲ�1����?�陇,S�heh��#IT���t��9�u��*y����J��ty®��4�"a�"�8�1q����ĝ�7m�vlK�o�������<��  �0���Yx�� 4�@�{�����m��&�u�2������A�­yB���&��Lk\M9�[K$�r&�D������9u�����H�X�5�]�u�¥�B����R���uD�4�TDy��k5��[P��D��{g�*'�)z��nM���RQ/q�Z'o�2O��]��QS�+}*4�FW��}S�uc^}�i����w�<��otz��ꮕ�I�x���}7��|�򬏑'�p��׺.���*�1hQ�S+���Qze��?�J����G�O�ed'�S�	�6.����ne�?�oZ��5(���'|��_�Ǻ�4'��J��ON�cI��cd������w�!Иy�aw��8�6�':'^�"�dͣo�G�w����P� �-&#N�@@)�������@ڱ�{��n#-Z�~��}\��#t�#��,���4��@~,��* G ���/���z/���oP��d,'T���I+
e�r��%�Ԏ���]�J�x��T�&]E0�>���ضD�_Y��:�Ӄ���� [m2:�tl�	�Ε�qQ�#�}��ɴ$�~867��I�4�vz����| b� �4�ᮯ�+�CIJ�%\��?��P|>J3O�̞�%�	�����Ig���t =�t��
\ Ũ9��l�9g�I~��_��;�b�Ο fE&l{�t+���$:2����� /衒OV��CEĮ��i�a�&�4e��V�4��[4RgmI&Cj�-h�mؽ4�f�������䗢��LyJ�|�-I44?���^�����wXl�a��_������ٸ*l}�~>��Nr�>�q�B�aO#Q{D�