XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����(���qn���lSҤ�&��?8�(L�ݿz��ijΝշxιi��I�ͷ@	�t;=�ƾ��A�������U�R��l�p>���8=��y͙*c4��/HP��.CTӑ�*���'�A��׬�?!�ѳ�4bh�����9T^LRw�޵�=�c��ng�br٥����Nu-�@I���k��b�D��D_��3�;����X�-���J�+6��L�U�н���U�Yƣ�3�A
���t�����]�E�.x����G���d�������˞�4@���J��5�t�k������&3ȫ)���&4F���_NO*R!
���I��3��kdK4عRU��u��bl�gG�L\�n�zc��gw�r�O�����p�9�լ��Ԕ��)(1��Aƽ�8�N����	�xT]��T���	/���#����.-�j���B����(�rDb�9��ޱ�Q�u�? ���Q��.�w��U��P�1��t���2s3=���s����ƯS�o��\�7YuU�e����d�f���Ka�?W����[�҃y�a:ɺ�Rܳ�f��5�'VM� �0;��b$�Q���޿��9Y�3��e��}[��Q�ވ/�H�=@z�2���x��\J��&��7�m��w�RV(d� .g�d&%]ME�lIꂭ%2%d�&��e �R�@E(�m�`���Ű�2����L�a�y��J��	?�����$��t'[gO.-��g��?/ɯ^N�XlxVHYEB    162c     8502c���g�`R$��J��S����沣����o�]�-n��i��A�&é�]���T���Vq睚h	��`��/�L�43��Lv����
�F�G�c�utw�W��̃�S��@����'(w��2���uX�IEv0 �Ax՜��"�)�;»7��Ǣ��;���Ap��6�V�B�\Lr�1:����|����r�)~pi�~�bFp���3cY(~��/����6���^9�Wu~y-.`��z$��-��NN��j��6����TD]���G�1Cm��S��������-hZ��P����B���p������> ���H�o)O�]@'8U�,xS]�s������O9j��@��-=��j�ȋv�Y���C��ߖ�?�\\,�o��ŭԎ�+��ZL�[p�a >��ig�*J����91К�b��j��*nբ�VgZ���Yk��D�	(�ۧw����7�o5=�d��&�l�۔X��7��H�g���_D�߷�/���|/ڛR:�V�������M:��)ϥOqU���� <�"���,A��$�+O�H�N��bǨ�?�HTޚ��յkl ��E �L���2V�IW��.��u <P�
u�c���p�PҨ/|_Ĳx^=��Q�ˌs�������Ÿ����h-�P��
[|�[7��Z�yA8q� �˨�xVg����jW3�CayOn�b�v9^�1�0��
�bu��\��HG[�o�?x���	
G�)��S��[�LyXa�u]�����e�����{�f�`n�߸kw��ZvfSe�����X�oQ��&4A*��$D��$G�W#]2Ɲ�*��D������U�͹��n��>�a���@�OYv��W(�΂e������FF�s�dW��%E�o�#��sî� ,~�fX�'c��8����9��c�w<5*&��LN�ԉ(Ƭ4��&Z�Vt��̢O��6�Iˁ��(����&����,NAM)Uq�-T���X�J؛�ZȜ���d�ݲ���@ۨ#])_�Rޗ ��	��$_�i$��d>��$�>��	n+z�\�[�����k(�zz1v��74T�c�Z=�y�/i��\�t�h��rd���I�L��]Nȅ,Mc�U�>�}����dU'b*���ڴLz��f0X+�;�>�z6�B��	nԿ���f�þ���*�'��qӓe".��Z*&O�=Rh:�/���w�ӧ5~� �$`خ�d�/�T�(�� �����'�)���O/�R�J�+>�M7u3$��0J����@���m/�y�
��Npj=��7��k��n8�婄��Os��Z��ŭ�j�K,<��L��=�7C�#Z���I����#*'?:����7�OY��b�Up�#�i3Bѭ���je�>��>%��^�sdB+6;5Fy��b�ӗ"��6����(���IrM�M��Rܯ.ڋi�n�%��c��s�^�:�DS+_J��ٞ�.D��/��n��x�}�7����͖�]�#i�S.�9��)��Ja+���qg/���W�淉�p7�~z݉Z��p����&&�2"�t��M?���G�^�߶��� �8�n��`�%�M.�����u����y�����`�Ătuc�K�`�M�eM��� l-_�I�~�DDW������휃��S��@��P>��9��Q��+Ԭ*�k�	�|��n�J.�&_�}%�n� ���)P�	���8���Z�l#p���-�*�h�fB��%_��@�D�9n�}Q���3��Q:�ק�+Ȏ���n�L'UY)�B0�y]�]��{T��p4 tt\�"Rw_��b���i�n�n�c�'9���&�&�Hn�j��y88+��p�Ax�b��{���;�3���4�u�6@�
Ee�6���>іR�s>��~D�=�k�*x�Ti�y� �7������)��[v\壴�Z�n�q���z��t6��_��j�u�-�T��8�H��u��Ǳ/�[�~�G|��A�U�Il������A���?��6�o�ۤ��ѧJ'�OM�~q��'+7���dy'���5��j�wR�}��r{����"���kF��E��