XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������Z�����f �� ������3�=y�%? �+��袧��qv'T,	��'�ä$���t<Ҿ�KhPof[~�+�z�JN��v�ӹٰ�E,8�+��W_������1�$Q�V�+{���u4<hS��#ڃ�R1�TKx*�MR�c񛾿����K(��N�͙��<���H�Z��iN�Q��CX^s����e8wN�N-�]�����k����$B\�����2'�L��S.ݱa�0ͤn�]��8��H\�Z�o�DI��u�A_��ؔ35��*_�� �D��X�D��?-j��G
|��ÿwac�H����6$�)��Q��F���ϋy+wj��Q�5?m�r�6W�7�G�
��N��=��X�]e�s&�X�[�/���2�'�����4g2@�6����@�q�ϱ|���pgc�"�Fw�Ž�h �!{���DA L��1r��6E*G�
y��ݦ�cs���Ytp[�%�i=g�>b%e�{�;�c�^���+�]��J���D&��$<�K�� �sYyv�dK�I�����M�8�r����5�l"Cy0<v}�ڍz�7o�(Ԏ(
���V��E��o�0:�q��6)}f��
[8f�Oi��&��~�c�C] !s�e�;������1��t�y�P��"c̋0����i=����~��T��{�q&]smʟ����W(�Q��NsG(	��p��F3�Ia���D�$���m;� 8����B��)!��lv�ך#6���6͒���6�SL�J��sXlxVHYEB    9efe    1be0��#��0�E�`�U^IQ�0�i���:���װ�$�L���8N�X6֡�#ПJ5�NQ[����B�olv9Y/����qN P��
�����Q4\q���ܥ��)�Q����B�o�>xp�����;ޝ��K'}��i�[��l��d��tG����B����R���'��rL��q$��*&���#�X�V/g��$�e�aA��+\�%b��9 �6��2wΰ��_�gٜv��@V��������=�ԷWtˡ�q��W��LDR�Ǣ�j����P�0T㬹ig�P�f<^-S� �Yi>����r��~��k�Ƕc�X˝�2�9F�Ku����^���-�Fz9u	��0j^������e�W�!EZ����h�z�)�j�����h�u�?9�YEP��tJ�As
)���_����8�RoB��1���ͥ�۱̕�g8�4ƾV:T�2Z }�$|�L�o�a��uL?8p)��U���?��g��)�Z(�s&�;�<Ӂj��j����v��F9��2�i<�z�w�&���8P�{~f�MNʳgq2��<k�)�ުeY
J@����ܶTР�H�ېq3�=Χ�ϼ��W_X4�6�:�dxˏ����Q�Eۭ�-��.}�V*��<_΃�T���>0������lW5�
���w�	M��%�`�SC���A�}�촟�f�yWE�"x@�i�0��ȼǜ�?8�S���.W Io�|d�y�st�����6�(����-u2��rٝ%�+B-�������95�.�X�fu��V�^�0�Y�kL�g�?W`�<MXf� �2 �,��vAS�kR�U���1�+=HO���ukn[k�����H&���`�#�#�9��s}Oq��k������7B'�����?8⡐ξ����[;��7}E_�͉�/$}���D�H{�v��p�Y
t@h ��~��CZ���-�|�|�k�8�hr��8���|K`���9_?R�kJ������2W�Qԫ�5r��ඇ����o��Qv�]�
B�=p'�0�dY�0/��'7\`G=u�&�9��F��/ �{�V6�¸.���d��	|A=y��f~���۳�Έ@�����^%v��s���
�)�}p�"�c
��FǙ�
�zdq�9�7��K�v����D�ZW����Q�6w$��O��' �8�H����%5	�$Ry�u��������ئ�؆��6`���L?0+=.g0\V�eon%G��L�hwy��Lj[���h|o͍xe��k�.12N&�
�61̦�UI�B��Skx�\J�1"�k(�����0ڲ�C���~���R)h�V� �l��Y��[!�HP{:��|;O��>G�݈R����$�ej�v��Y���(Į�8x��.�m���3g��I�2����wX$�N;^���Z&���mA��
��y���#u����扤��F��5�qR�Y�\��c� y��h}K)���0�{V��؟���^��ucE�ǜ�!�\yx��]sGOc5�i��ۅ��
�a b�j����"��?ǷM�I��,���=c�O���<-�K]㊲l�>�Xc�k�j�f�������A:b��&���ٽ��}l��<GG(��&��+
\W߶�T��y�ƩW���ݟ~���`����)����.�e��������d.;���~���$j�wpn�r '"��d��f�2s-HBO�����[���G�S��'�;-m	���B��9��&o�7��I�@��!�n��P��^܍e�b�(�i�Jd`��=Q��c��}WOH�i�)ڷv+�X��_ޘb(��$��h)gȉ�ƮYfv4�r���gk��?���iG����UkH�9����מ�#JEä�f�N�@z�q����ȑ�f�|��3�͕�5a��׊j�5�=V~O:����}����JpF�� ��K�c,�Ĭ_2D���3��Q��M�Ds���:���9�����I38���HG ��fU�ܨ�%(�����k�Ƥ�S�����v�-r�@5�O���|[�򛜽�V�����9_mdl7\XL����QGAXj�Q

GC�O��>?�j����p���ٙK` �����q�,�d���H=��"���#��F]lU�4�{v�n��ʾ����{�YdbR�za���,�b�ҵv��0��\hn�H���6�<ÎXsK��خ�陣�`���拜�uP�]&�q�C��}����W[s���;_��@����3�h��M��i�T4����/�DX����]���듚��<ݜ��QX�Bï3�ʂ}0"��a0p��iMS�ۙ���<��� � ڛQY�0�q~�V�	(L-Pv�ޙ���(�|���V?������^���I�	�A�;a��Q�� y�	Y&�g�É�b����!j\4g��CH�N�l�؇+ �����mG��=?�x�=ޥ�����\�pbQ�Kͭ�s
|��+�=��}+����E9zTe���y�$F�����udf*Z�k�*aL6�ި�b^�<��h�k�l/Z�+�/g�2��Kpxg��.������JiI���=��ƻ{\Q|IKn�h:]��bz!֧qJN�{Y)8eY(���{8�$U���@��r�k@�+��+[��wL]�R�� �C�L�t���2*�����(��eE_rL�(���"�r2�A���N�SB;.>� �c�BzD��}��2�'�)!�KƟ񼐲���E�h�g��c��NL��J�HK�Q��pU����#*W����'d�
��5�VY!]�;�7Qj��n�*� s���܀3n�A	�TJ�M��.|��b7�r L���e��%����tڱ��+�Kw��\��9�2�h�m����?�GL]YK��9ہ �|�he-�2�R�Y3�-���u�0o!%T�h�ʼ~�FP�!�4�&�
�\�;��\Y�̔����Q���xqE��e#�?Ιg0�4U�Q�ԟQ��$���~���T��jI
$�k�A����#0���s^Qy�+�����g�MÀ�;] �[_o����,�)��@�'��y<�r�mq�He�2w�
�Eޮ�}�)ߢ�����L‸�$�u�"��\��q��m��@���s���Sf��|Ա��@똭(<����I��7<&�P�!�EH���1���9i:q-���-�4� 
��z	�L�R���Ǧ~���,Cm���s�U��(4�����CGr��!]!����}��;�Dl�ϙ�]��g��߹�2�ݡ�?{���q���"sY^_���p
D���E5	a�z��X5II=L.Ѩ�hpӍ���*H�~iŖD ��@S�y�m�Yv���uD00(��=٩9�z�@˷U��o=�O��Z�� �'+�X��4<L��z���QkJV��`+O(���$���N�-�x������p;ҿA��O
��3\�A�+�k��a�j�%J����+F��B�����E��Bj'�7��������_ح�/�#��~hI��9Wf����T��W�,�Y�����	'�-f~�D;��~��Q��d�%�F!������m�J�|�׭�SMD���� ��j�UWZvYfZ!-�����t�c
���8O�KR���V��F��|�iO�%���[1ے俹�\���:��@��rC��A�4�o�#����K�º9������b�����<��rcgf/!蛘ޚGE��<ںH���)W�0���I��q�w��%k�+�E8�ѽD��8��{�I�K)	���D�fC+�?��Ӣ�@h»[h�Ro%�"J�7

��<�3�ڐfb,��q��XΌ[�%���Y����Aţ�����2��91�M^�Þ�D�����u#���
��bM�T�Da�%q��#�^�F��C@�Uy�E�`v62�oxy+h������~W�?��o�1`��f=�v>n��"�Z�7�0���~�.���а�˛�s�Y~�w�Q�%!�(��kq����@�XD8&&Ch������=Q�}���=�v)
��ߦ(9�E3���^�6F(�7����Eg8NRb�靑"�MZ7��9��6 �����*C�;�Bx�1��i	Q��L���{���<��ڦ��2���VA{��nZ�M;=��X���\s9	}�GNe����|�׌҂�<_L�'���CHS ����ؠߩ��6����X	�&� q҅� ���N�D ��#(XH��|�<jG�p��G�P�9��4�:d� ���_�~�����l��`0�����㍆q�wM�G�>��a���M�l��j�}��CDu�G�k���-qh0Wy[��r	�Y�إξ���  j�QI��6�?,�*�Ll"��[踟NIj��m���,u�F�} ��8���1�Ci����L����P�ve-ӿ�S@�|�H^_�A	:Y��G�+[ϟK� ��|��n�5$�TQ2�.�Iø��0շ>h��b��H(K�W��m��e������8q�mv���F�m>&�
*�]<���2�"<ɩҵ��u�K��G_a��T4u�*|�>p���[ɪ�`�+�9@�l���6@>���Y�C��P��i������9I?!�"7	G�V��|�D�|���Lݚ�1��""�숒���2�1�>�WC6�}.6b֓`Ŝ�1��
x�D�>隹회jS�q�'���xZ���W��L�3FZ��tu��>ǝqdz?x�V��VB}s�1��:�/���.T���Ǭ�H�,N����<ɦ�M����"�.@��N�\>��a�O�^��T��f�U6�o/�!e��\xʳiy5�J���82Ef��xc���O��H����=P��y�j����F2KbQ�ԯ|�Zݪ;�nG1��u���T=n�J� ���i3nޫ'Zv�n�1&�:�K��:�Y����0���r��L�#�o�S�/�n.�%�6#�gh�#����/�'Zl{���~%��'ɜ�N��B�����S���E(����Qk���S=�J#���͢4�Kg�c����)`�	]H�|#��~e�,�|k���@kM��cs ��4�Y��,��ϲȉ�L���d�ѝ��?�p|0%���[[ǲK�R,<��hW5�cj��O꫽m��bʣ�]��)T�����9ۚ�P� NUl�����%9+c�ۆ|���(����|�߆Z�=�Tr&���{.�Ł�_�HzX"����.jg�1_=KK1�i�TT�F=�2������r�(ǽ6�u�^�g)�����3��'a}��6zZ�e*�x�����v���6���H�V�XȜĴ�-d3���ʬv�Jq���KN!�Ϟ����p��8�үh�M�sp���4�ҒX���S-�g&�3u�˽�M��y;	8)�4om�OI���T{���Q�eL���8t��o �X�^YJ;����&+Nތ ȜF��	>��&Y�I�6壎�1N=ֻZ*�H��G k�mk�~�H�/�y4}��ïg�ɤ73�����%8��`��>z��?�֔�!� Xt�Ý�.}��C£�����@�w���B���Zy�q;Y/_������'D�#833J������I{�eD��{N��x�ō�l=�n�]��-��j�QI���/�����]�%����Ȩ�o�kSm C�O��0�f�߳�u�n�FwU�����rc�	�Q�`�u��C����JR� t�N���'3�=,���	 G�5/�
K(N�!�X)�]�=��o4���ОG��B�A ́�l���rWc�a|B��hz��^=}���H�C����jX,O8ܽ�������f���k|�'|!�-�0�?�X�9Lh����xw�,=zJʖ��S����@`���xa��R,���+�(�V�^�h����rnq����hL_4q���kax� *��^�������wP��g+�j�7�b'9~�+�����ѝCzQ	���'��/�x{e���͍�4~���D�=(*|�� �(�>��;sղ�-$B�<FW)z]����h��W*�H[��su�&��Ώ�x���� �.0$�F���7���"�؍̺~�Du�b��7EGr����A{�)ǷLL��_�̕�F�p��=#+�q%��@$\1½8/�;εo�����_#�Ksb�y%&��c��f�{�^RgW�]�b��]�`es��a]k��N�)_�|=u��r�HYO ��㕫�)��ŞE�M��o,3���d�`e���mc��F3`c3=���?�M4[�В^.ݨ[�/4b�*�"#�@����L�b1��k@�*��>�;�.C��s��ن����_B�y�1Ea���=�=<Oҽ�́Bf`�������]QP�X�P�A���^�|��H�,dx)��9����.���6���5�J��<ٙD���I)�>�Dz0Ŧ��jVb.6�xگ52�n�g'�_|Z��Z��N"�1�s�um��P燥�g��.񞙄�,�,j!���>}��3�����&����ҹs��G�"�.���Y�x�Tn���X/:�70�$F���E�;S�I�h����F̠]�k���
yBE��Y`������J�����Z����oh�L�!����lY������`n~�"΢�b`9�;�O��7����q>���p��%�Z���J��5��م�E%����M��n��|�h����o��k+�3�s�εo�PK�h1n�D��X;ȫ40m�8�U��Sl^v���T%iM(=}�ع���fm�󕒖�2�a�v��Kby�?A"�0��oiP���Y��I��o�X��A�F4��mvq�Gx]w��>.H�-I�9^�3��ed9jB/+d�
�Ar��K�J�t�Oݟ�s�6D@;�Ǥ�W2��xG'�nvⶉ�s?y�!`��h�I���':��7{�T|v�t�	��V�E�$���Kd��c��߆��]�m����>���Z���\�mDi�8���