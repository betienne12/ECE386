XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �.K��� ��_-d��s���e�O��%����U4�3�!�1S�i2Q�a�a�a:Η?�+(ϛ�5=z��g�A���oK�&��ݓ�uձ��L�͖��Scha1�
Z����=G��
�[|�/��n�-_��[{��@���K����ˑ묕F�pf��)���ܜZ�Hz$�Y,dFEn�O�fc�S(�:��Q��jӐ=�<䳆g�ŕ�W�Y`�qb�5����C���\u�G��둰����T�_�-6��r��
%��B�ԃ@R~���P�S�	�B�I��5�VFD/�$�$Y9L-2^�E����M��A���ؿR���ДTw���Ϛ�K܎r+!v�2c�; ��H��)ؠ�i��#�971f:Lz�����s��։�c2m%����е�u|L��^w�iW�a��%��2�T_����!�g��G1Ɓۍ.�?����,a�	m�L�h77io�7䤭=LHԾoK���˦:���[7$�V�l��I)�Ut'Ù���	P�ԑ �݈6���A*�����*�Y�����G���*֙g��-N��C�rXb����׸o�V�J�T���p��S�k�&�怩�(ː��-�6�l�B��BE.#�ws�X�I�.|5���Ѵ�j�ݗ�i!����%};�e0��+ѽ�A9S��[�w�~��s"4V]@�83h��M�:e_}�̷GP�#Y�a>G�|:�	
8�>�{qT���.c�Ç��rp� ��>{]��F2��1�IgR;��DI��XlxVHYEB    fa00    1fd0�~��<��$�p���h�؋x7:�U >@)z� ��)d�(1x|K26�'e�V�4UI~׭)���%c��9-��f:�@ꃫ3	�]�6�����8�GW�h��'��L`DEr��~��1���*�-&@J7�Q���e�IU��]|34�~�.z�<��P��r�?�����6���2�c5�is�q���J�?�O�!|�+q�B;d��|S�d��{I�`0W�H��ƕ#��J&�Wc��טsu[O��������I��Z�W���+,LMKSPUp�l˒�A������d^ؾ9h��ѳ_��¢'[�f�E> B����ɟ�^��I�����HT��p��3Ԩ�#��j���m$��b�� !]��ۀW�V>�-������K~H��$@��.��X�X��u<A+����(��e�q��4X5C�����?�ٚ�=����I�aխ
י�����lp��4�-\Ry� ��ȷ��as%���nT m�����5 �`� �t�w��ؕ�WX��J|�E[��U�R��c��,����]���4�Yxc������4p�ا&J	�!���oh<!��{���t��Lq�J��N�vF��28<o`��m)����2u<t������5cS�zjY��%���᛽�D���%�3p���5t�O��@��Fa�Ն<�����щ\#���;��������_�ѐ�����;�=�.�f�����f�1���":h��P��,�֡c�&�LR�j�SQ�������E5��s��GC��"�	�O�Kis��v��@���գ4���e�X��s�ګ<}i,��I��o��2؛���4����V�\7���Xz�4���@�����l���*v��������7��gs�H��<�����I��TZ �E��e � n���^��O�6N��'�� Z®�E;�lM��;��%[�=9[� ��e��AK�]ctb�dfV�^q��ӑi��wh��y���Ꮵ�w���(�KX��� Y�K|V�m���^ ��0+{%>��%�/�}^�&z��ϝ�t@3���n���cC�RB�[�X"�@�ȀX�zK�y�X�F�!��l��W� ���~b/�R�9,�9�����p@֊�h��bJ���&%�!��7��]ra�?��b��~�_�����2ݕ�G�|;�3Z�I��\l�d��h��ڦ?����vҪэ���� ���]��f�c�j6�����!�����J�ee����7V������Q������Bp�<�?n�*�_�/L����iQ�PW����<��`����}Dڅ�FJ���^���bQ(�6kx%5��?ӆ�!���ɔY��n�c1I���M�E�r���_�	L�yXVǵ���
w��~2/٧�0�B�&xZ8�V4D����A����iN\b�Bݑ˲�$�"ڡ� �A���{tȪmc�`��75r]U�"��*W���E�	u��=rɫJ�_XqX�Ti�������2��w�&��H����ф�ЈP��G�ӄ[�e��8�Ł�l���T�o)D��M����Րh��o�`(Y^xȓ��"GB�?Yך�y��1�w�/�/c�YK2�*�IE�we\�Q�c�����G[��kB�˺�2�X���ח����ב�KLA��r2�&.�F���H��:���t�H�s��hW��0�����{'�F�S��ޒK�
�
��7�@�	%���ib4)z�M���
�.����nbo�B��$��эƿ�9e:�-=�NV����Z߮'HQ�g�|�U���I�z]�{^UqU��l�>���3s}4z�.(8�ӄ8�'�E�(6�N҈Z�
�'�?ЁR����+?���Hl�D�=�+z�D���0!ON4�0ģ�Fg��4����62���g����p�t<^!#GV��A��kP�����',9�����d�3�F2\�	A3�饂Ӝ�&��iMoF�J"D�!��ץ���^=�T����6�С�w7�{D3"�hN��Oz=���m��޳������h��Ɛx�t�p�.n��[qӫ0ʨ��!�n+�T���Gl}dGbO�|���T��$��?f�Ζt<��q@�>�a�F�`4礵�Hn/Ȫ�2|S���n8�2J<��4[M�#��� ��@�r��ӏB��LDjԐ�9�V�?%71� �/��&Ћ13��@�	p`tK����{$�Z�E��V�1�7 �m���<�	S��fu�{\�j3 n�ޏs�P��o2�B��f��}�#! 9�Zܾp��H�����oR����Fۿ;.�����z�є�Ď�	:��������y�y�rI��R����&�t s���Rv�*��E�H�bA�ϴv�V��IB�7kN�����	��4�$v
��'�+����,�N�4�@7��JBƀQ���5�Y���.�Q\���+?
yÔg<̅��7UU������=���n�t~>���}I�
��b_�W�"g�v�"k����e���V|��,~��P2���U��!/6BlmJ��(�E!}�]Sơ�փ(f�>0W��ϧ�>���}+/S���Rv�&��~ؚ-ߊ�&h����#s%@��r\��S��.���y
 ��4�꿌|�w��ɰ�IGd�������n�0�NkL='=�!Iϟ�S����خ! ��{) ߌ���#';mK��;l���o.�칾Jc���O��CV,F9��>d#�71��Ř+9�n^ؽ1S��(�t1���h�O(ȭ��T��3����@��D!�\U�͈��:W%�B�jjI�؞���qܣn�t�y&v�.To�#F�uz�!K���Q���:L�$�c��s�}�!$?7I���ͽ�q�uyK�,+%�]�4J,��b�ݢ��]�^ �m|�U��ƵԱ](ƿN�̆y�Lzn���4�X�-%!(@����X��j���9��6�9�h��x�s$��^���T��WWK ��1���A� g�L`�"#Q��H�\#�����&b��r���>/�ӟYu#o$D�J}hO�n����r����%$��o�R�q��[.�o�����0Ԅ�|>0�k��_�CӋ3�q�ni��`1��	L��<���������.���]���P����,����L�_��M�K����{�)\�,�H6�" A��G��&��C:� �CoJ�:n��j~�j��;-��G8���`=��/���ٺ�+�.o	f2�͝�M�������Ǖ.0���c�uN��K2�P~��)Z���ơ��i�J�������h�^�y;j8lѢ����.p��������X�N��j$'���_q�����d��Ó�#yF���x�Nq��N��,y\A�����M�[:��z�TL���A ���7��e�u3�\�iXՇ|/D1-��w,0��$B�LF�=力��y(>�|4�����az��G�w�e�I��Mg���B��GS��=Y�l�u��K6��i1}v��F����a��?7[��O꨺r�������ދk6	��?��D�-`��]���ֺ�P�U�@���{���h���6����I�AYJgkjӥ
�%��񲩢�+"#�u���6�c5ߑ6AD����e���q)��W:?B_����eS��ח]�9)ewP��Zĩ�HK��)-ӹ��3	�C���P����X��`���,|A���Ol�3��B��n�s�'^&C4���'7|<vO��z��>9<I���C�D��i�����i�2Q>+���Q�lM� ����PDR/u�>�~�഑�q�0�f�K�΢�@���^<�<*����p�|�Ȅ��/y^�G�����K:>����X'Snzmt���������vɼ�3�pĔj_���/�n��3��si����]��Z�Is� 30o��=n������"bh��TX�Ƚi�/aHt�f�J��q���C�a���7&�l�*�����๲�$�]�J����U���@.�'m������D*{GN��X8����C�����������M��X]S�7|49f�^ �p~#f���<�U麳Ҁ�����Pw��Tk�Śog��tt���׮D��rE?��J�A<g����+B-ȗF�X��D�?�N�C�Cz玑qTMS�W�4Do�5�zW�C��R~ә����z��@����:�i[�ʘ���#ʚ���W!!��l�b߇�)�2[�1�՛�G�������}����&ϟo�.]yz���_��[%r��W�I�a/bD��!<������p��l���O�P]w���MG�lA1���po�Xྑ���Z
j�:pV��ϝ.R찘1������*�&Y�[�Ԡ��>3�^0m.��H��_�}6F�9�m�
Ϥ���0�,��A��r��q~�`��H�.ԋ�s�@/��n�l�w��Z�;<�}��9&��-���A,�؅B��������;�����vof��%�Y������5��T0�aY�����R�{r��>������M�z�_�j`�1^���3�L���gO�U���(1h���p�/����=�"藏Kg�»� ��%N ��{<�6��$ܶ�¾��}Zi6y��݉��V����OM=�������%��,5ш��/�zsQ��b?����<w�T^i9�j��V�;����^�S߉����qޘH���!��:yC˓�ؿ�.���q�*�(��-w�������^��;�=��y&չTu�oH�,d;�N�)��5D[ ��f<: X����α~�|/"Z�>{�D���Hn��eߺo>.2c1E�iT�O"���Y���7�؂2��9�^.�v#z;��	ۏ�pZ�7�Q�b_��0�c�|��`�Ĩen*p�s��6+Z�l��O���e�+6�C��)�^�a$�����n����Qd�n�zF�P�甚n%��r��o����&��L9��:�O;�`nЬ���N�ۏL�Y��&9Ê��w���3�Z�V��BZL�D&�<�5�����_J=��hx�d�Fh�H��X6
3�~�I��f���Y��5����۹" Y�ޤ0�Q�#FSt
 j�'D���4o�A�8�Y��
����P���]�l��rN�Υṥ$�w���y���ia�x����+}�W0�4�V� $�������xŗ��L��J���f܀��0��7����Q*F��j��}�-������L͗�p�Q
`�6҄O�>s}ĝ��W�!ޫ�����dV�Y���j�8��� 3'{�J�/�$c@���$7H��~Wۤ�L�	�#	1=k���^1�_�'m�	�6Tb�T����ܩA���e���<�AG0��rH��o3YK�����x��;��˫��k��I&�K� ��6�<�0�A�!��G��DY$��-k`e>&�:����;|�ޕ>c+���>Lz>uW��tK&��b������O�Lytwn����Y�r�EU�8�����z�X��h�����k)��C��_~��'rr�g��9�̞�:�E-��>�(i�] ��QRq�%a�,a�X��\��*�@>k9��R�y�Pc�<%z������y{ڨ&:�(51/�}����q��/�Y\G��R�@%��w.*��
��b�Xٍ�iĄ����c_H�����i+#�fk���}�����pSN(���R��Ж1�NJ���n>u��A�c1"&��ڋ���7��ʾ�+��wx�o�M����>^��R����p���[�l��8_�su'{6��1VA�ՕJ�a/��g�;�/���*<��_+�'U������svJ74-k@�HUf���k_��h�T�7�x�Z��4R�����\W��M��Ű�5�U;W!��z5G@����o�Glط���N�I�I�~�?�nbwo�2K.d-�3n�1Lj	���Ԧ>��Y�����ם���,bj�W� �I���e "N��<����/gP�ڨJ�J):II���5��Bp��8���g]�� qƉE�2"�67=}�Kňī`��j��������Ov��ߝ��8m�Ҋǰχ��%�V�2U��D��.R	�P*I#��)A�t>X��R�M�9�P�0O~c2�5�y��RMXܜ���Vݘk��Ԭ�� �8�,�6��]�~� 9���(�Eu
�g˂8�e�t�Ͼ�*�v�}�|}(�����N\����^]�m���[��L�x�4,��	�I6"�|��5$���������P�q�<�M�{$�%�$����ϗO�5���)VE�5�x�j�2�ns���/a�;8a%�U�|���}����|P1�c���,OX��JH�=U�g�W�Y;-�U�! 
���s���E+����p1�BMU�в�|8G�������gJ��>G��U�g���X��jp��Lr[Pފ���1)`7����oRՓV��Q�c�n�mJIe2Uܶʯ��J'm1��0�R�>v�mc�!��M gX��{l|��'S*u1.��UI�Լ#���~ijp�}N�qK;�A}�4�D�Ad W�3O�����	D@�|4ߞl���!�0�.J-��3�ə;ܣ0�����\��n\�F���KF�Z��'ϱ�I`hҶX��y����@��>-M\Ԁ�<w}&8�K]�̅�V�~�Ecco��;x�M�XG�ݨl!L����!i�A2��� ]��i�R83�ݼ�h��dG��+�~#s��;X����$(�Ie le�dR�߄T�=9��Z�!� =z3{�غg��{-�X+�!�[.�&�\��;MY��t�'����kP�4]>f�3������"뾲��s�d��y��n�m���' �v����$��ei/6��]����Xx{�%$ra��ӛj"��kD�o���k#g�Uu�Q��Zϗ����rQ�٦w�G'�ëi\����ـAb���#L��n*��d�m
�vݠ�L#�/�^ݶ���+Vā��	��W��r��&��&oK�����S"�u�Ʃ�;�d-�m�)�2*�
�Kw^�p��rӫ �ʷ|���d��Wq�zY�
`q�\�q�X޷"��d,:���>�qk28����-�\�����V�4zy-Q���t��.�=�͘���j��C�����0 ��d<r�K/%=�{'C�C�};��7� ��4�RR��&.�:��i�A�(��p�_k$r4}��hQd+]��2���:'6#��h�YA�bQh�|7�����C�{L"��%�G��e��Ch�R�^�[j�U�1�'� Q��/�J��x��Ce&y��aSl����j�4�Cò��Ъ E��5;s��)��N� ���lT̰�C`����z�.�7L?.Pаv���5� �W4��r�F�|��GG����0L��t1�J�骸�P�}VzΥzEM�!jWhk�T�<j�6�ZX�d�:b�2h��:�c�̶T^^���i���88SϚ0V1���&4mY�����g�UR�5Z8��F��?��!a
�/a�=G~�y�0id������֧-��.�o�o����t����G!�<4�T�z�v�9-@q���}����|N�2*z�$�
GY�n힚ȁ�h�j���%�ۅ_%���z�:��)��`_�=�le-\i6��
����E�L�!a:����Y܆R�	|)�W� � 3+{ҕmŊS�{[��;[I�h�Bհ�sЋ���Џe�g�E@�x�)��g��C�	��"NI��%���_��%r���ss�j|���g�[y}�CHR�b
%�Hަ���}*.�W^��=�.��ص���?/�d瑆����?����d[:O.%�b7�N3wn��PN���9��P��S����6�yk{g|��Q8�Ə,��>����K�__�P���U�̰�
��b��{F�����^�*����x1ez���M5ן��&���L1�aFF�!H臧��fz�����+�l��
v{��&�&o�}GBD���H^gM���Ӆ�+83q`���D��0�%���}�Z>/:�'�zXlxVHYEB    fa00    1340w��:"�Frth��!�*���>�Ո�R��$+��nS
�:��s�ЫY_���bI���V2{�.w���N��k����^G�#ܽp��3�o^�F^��3�Tc��do���D�:�9T��q��ܿ�.�/�wOÿ���U�v��@���Vz4p��P�J���h؋u��Ɨ j�}�p��^�s>�H�_��Y�]���}F�G�5�uDpk}� bؐ�eAJD��d�|.�[��F��p �D3$`�,*<�u�l��%�o
,j�}-��F�9�P��a�����H;�rBҌ ��y��^��)��F:+ʡ�~��]|���I�L�Q�<Ez|���F�e��y�	��݉�al�F:���x�����Z���G%�]zt�)�A�}�]bZ*��E�vw?P�K��J!�ø�S;�::��e�J'
~�܋��o
]XQ�4�Ms�����d`s	�0��ƾ���1}").��]�{A��b��U˰�YO�(�+�(�OX)\��6����m�2s*�2�ORφ�Ͱ���M@�gQ��.��U���"�wۡщL�G�L�1pթ��E���P=�P�!2��*�=د�<�`��i�Y��8yU�?�t���x��E��[E�`�]D֫��k-!����y�����>�^D{�Ws���mg��s��c�z}/a����	�:Ly$�� 4�+Y����w���B��y3rok�~�]f���TB`��?�NKsn�0l[��]��c�%���ŀ��T9WU8u��+���Q7a�&�q8�߈ �﨔�/Z�>b���6����0�l�����IMĢ�5�RyUe��a;=��4L  l(�A���孆�5dD����s<����q_����cƢ�/)am�g�����f�:�t�ϕ���"`�3��m;�m��S�0XZW���p�R͏��j�:��|P�ׇ��8��l��;��D81:R.����eK��㣾
H�H=cB�6�Xq����M��NOm�1�#őH�#�Г	& =���E�趹05'��� �w�3үqFψie��N��J�|�)��� E�1
�p^��=1�_`�4��Շ�8��Y[p��z;%7�ECCV������(X}�ЛI���a�[�0�8k?wa	�[�����Pi���G��ˤ�VF���cR��G~���S{�]Kw�,�� w<w�\�cK�MY��E-�r� �r>�v�?�?������\��NwK����Նqm"=ÌX�!���^hQ�7�GO۟��M���Eh�Q������4��ʊQ��U(�O�8C��ap���ŻNΥ��w���QKo����T���+���|�qr��|��י���-�N��ɕ-�����&a� '��>=ZZ8��%z�'��d	c�w���|��0�Q}\	��C������!��w�
/n��lc7�����<��>��Q~6"�x=�?�(�)q�֭Y�hH����0��
��ZzR@	ֺXzS7 w���x�6���[�%�5��d���<��)��ߎ�O�p����B�cM�������+�����Y�O1.+�<PD����
@[C�Q|�P��Z�����!y����"� � ���@����i�
y\�u�NgV4�c��2�a��!�˼�q[v�p�U�q��hq4~v�B[ �݄g5���Ax�]�7�;3��zԵ������`���+%�"���c)�ˣ�`�.,>{��6�����eIՋ�գ����|�C��a�}n}2��rOn�Y�#��:�Z`]ȼ�l2�C))��U���k0��Էw�d�����<���uv��0��������޼��/t>vA�CzY)6k�-����ۧ��׍̓i�x��e��a��˕�|�ఆҼ�s�#vb,�*��Q�q�u��=j�Bާ,�A�m��y�',9𴔣�ʺzcS�������۞L[π,_@�g&������'�=�2l*6,��v���z�u!�a\�ޘ�ŐH˯!�8�7�F y�ɚUʉ�h�I��1Ρ��� �NN��	(0��ܐ���y}j
.�x���L��\���K����#�T�~'��ťE���F�R?<�a9��6�TzT� ����Ð�}��J9g�_l]3�N���ģ	�8��M�,׺��9 E90�Ⱦ z'�0eZ��,c	��u�mD�|b3��nҍ�ň��ρo?l��`c�tk���b�M��z�����
����c�4r��UG�P�K�,&Ul�X���Hz�h��;L����H��F��x��og~>R8���4��6�V�.���~t`��}��`����@��i��H�[�k)]�j;:h��!�%]��̸7�C�x�4����|�pf��޺Tm�&�d>���!J!��F��1�s�.���\m�S�m��D�M�ۀ4b�QN �5���R���H+��UQF�/��I���_.��I�Q3g���]�!�p�1���F�ϛ��-1	�ڹ�U).¦���'�J63��j�����Ap��>�P'�I������E��H���,;;�k��6��?�`4��]9�?�H(����'�+N����o(m!$j�\��$�1�T0_\����;P,����r\��'��E�a3���T���a���N{DI��$���绤W��hX{���.�@���?��h.�ly��y�E�z"���:*�m�Nj�絮PwZ�m�u���gH&�q�=�{_�d����6ܘ)Ǟ��X���'�Az���A��?�c ��6�O���%�/M�Q�/�^��L`�{�R�n�u�Pg1� >��1�7�3.��d�ڼ�L��<�����Л��0�����>�|nY�����H���0���B�D:��|�Ч��i[絶�� �oY�
,;״;��2�y����0k50���-O8H�RMw+1��a�·������J���e/o��_����O=�����c���,3ܞj���z���w��f�(5��h�*��Q�E]�i�8wUe`o��
(����ܬ�Y�2t*���I�
�P6Y3v.~E/��OM��[���ѧ�X��}*�T�����و-H�N��>u{&����cT�E�/�~sΌ]s)��틇N.�:Ƃ���SvY/��4�I��Ϙ�k;�|2W�ֺH�X�������e�vi��Tc(��Ć2��[s��4h?�)��/:[�p6��}�-[m�{���.o���$�%�`|fL�������eQ)�4�hqA#b��n�ļuy\ s���^����_6�����V@��៭lg5�?Z�)]�6M��B�H����ᢱ�֝��[L�u���G=�f8����d�n� �Ks�C;��;�d�&�b����|D�ܰ�{+�M���.�cB�v;j5Q�=f���?��H\!�u���1y������͙A�؜j�Z��R  �6�H6)�4ȉ�I!����F�J�Sx8�ΐuM��/���?�@���C��$>��e�6�
yfb�|��xn�?1�#�3�-K�CW�6�n�$�`D���UmϘɛv�w#2�ҵ���}�`�-�����k�(A�~Ω2,��q�1�!]���բm�� �b����6���%��
��+��(�����]�f4#28r"�7� =�HW��P�
h�F*�����H�Կb���	���Hz*ٸ�؞�sF`{�UW���y;�t|��)��PyW~v��z	$Zu�<�AA���ac�{�3&l�&ŷ[`� ;�5m`�\{��J�a�x���*gRs,A�=��Ů��n�i@q����^���R�YIRq��5��\�w�_b�����w��}��L����:�h����`pQ�~6�9�)�;�D���̳�2%)��O����},��rpg<ls��ʹc:qa�)���<�1���{C�V�ۑ*��g�k��Ջ �L�?�^Y)B�r�jh��VP���\T�l�R�����$O�<V,�B��]��6����� �����P��rA����s7ӄF'�r%�/�1��b��ǝ���$�d�*�ۚY�`�@g"ti����1X0s�E/�et�Br���(��f��>Ƞ{�S�r��I�]y����2�mW�y����/#�arnnD;hpf��sx��Oi��tL��%l ��E;�Q���'����n���|?U�A����sΤ�ּE��\�K�Чq<!3?f:�U�����8�[1^�����?����<g���`\@����ϘMp�,���
�o~HA����ܦe���V����v���%��4 {�Pݳݒ`d�������^E;N��y{�����@I�^� ��I�)���!��褥Y(����"����N'kR�#@��'��xo�S�0�L�޿/����
����2���˂��o�� �-V��}3��Dz1�I�յM�N�(I����D�X��<�ԛ\�b��x��d�q�C�V=Iaƾz�aG��$�EdY> �MYE	�Ԧ�j+	�t<N��*��2+,��y��թQ�!�+�����B��pH�X�f�j�0��=?]����b[a��ܙߦw�G�*��{��m��s�a#5g[��i�9fkmjDlfk�ȓݭ��d4�ẋ4�x���!�Vķ�r��ǳդ{O��vLq:q��%�GX"+3���WJDY��2�ǖ�%�7��c�7�k:����v��@�aK�6վ֜��vi=�(�?	�}�ϥ�(��F���%?U��a�D����z���nq-w�ڍ�A94���\9�eg�7��� �|�5h�W�*H~����Tr|�#Ot_Z�{h��p���fVf9M�q�w�O���<"XlxVHYEB      e7      a0J��XZ��K0��u�vm�p
�+u@?�����:\���_���څ`ux�A�}	��$�O���stsܻ�$��!�͖�׍�t�v�QJ1�;c�K��V,��p���v����C-�.�M��A�$��Ǳ�Vӵ+����k���A��H�!|A͒�R��z