XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����I���>B%�rPQ�qZxbH��v��:�5]z�C+�G,'���qn���[�|����@8�㾬f���_䏓NAu�)�fK�-Z����~�?%/#o7�K�U	m��)̖K�˗F�}�d����i��[~�f����\%���<}������)�Xn���?��ُ����'�)�giM��rQ'g�_�pn-�&��{TZ�U�z�����Ij��Ӿ��٨�_�\]{�]�~R󢮤%[wfΊU���R:!�(����~�Rܚ�>�Z�UY�ܜF߇�4t��@(���8��S5f+?f��8/�W`XB
���^�qn��َx��M�mI������Ta1c6����_��Zz�P�D/(ه��E"WvGw�U��Mѝ<C_v��a�f�����CT��e��:~��.�M�6_���ϻ�l�ɯ�Ad�z-����\����z`U����ؖ`�� �*���xi�����eq��|Zrp�Ę��;?m��YJ�ܶY�� X/���U�"	�]"H�	��Pm�ڃZ&�`F���"�.}�܀�rz=ʋǤ���"���%��,&&�h	�'sK,2Q�Xw��2C63Z&��in�s��a�j=VS�!�R��:�^��Py�� &����T����>��s�?/1z0�Xy�d���nC�ת絰���R#Pq�\�20`�ƍ�;
oxd�Db��������𹳫�����_��4z���Ƞ��}�2�A�&)�i!��ݽ��K�G���`�XlxVHYEB    fa00    1f80��~�د�!�=����W�jЉ�o�\���(Ea#���D�܃�5i�]�5�9BQt�(ݼ�Û�o�4���\�����@��']:���ᇹ+����2[]�F���2���'�q]�"R����i��@�M�zNQa�݉�õ?s��-��C^��ag�E����[L�F/ �tܕU}x�P<gE�wz����Y�!?��P�˕����$|�|�ĹT>���1��;J�~r�q%Nu?�f�e�n�m:HN����}\���� ���N$0����6�<�Qۼ���lo|/�g�&�]5����A �M��ؔ��֣#�t���F�CD'��F:�!�M���+B5J��4�D.�K���/��>�wAm����3I[��jA��\�;���p��-�I���?-�����V�q?�~��L�c�\N�p�~i�<~fG��s�}�Sjl-;��5d�ݜH3^"�T�A {��)�C��,����Ωq?���٧fp����>�V�=��ze)Ԭ�}^+ ��C{�~�=�;3i�Ȏ̿f��oF��c��i�`���KN�J��HL����V��G�>�4>ٞ�$���fDoP�M6�W��0m�K?pK�俛l��?F��N�B0b�ܒV�l�]�����Hw���O=��^���r��v����Z��x2lKk���Դ�U:Xx��M��]s��l���7���*;���f�nOd2��'Ij�k�mﰑ;'(tr����w�tQKe�W�����o=e��9���/)c�3��Q���Y�Lmm�zg5��'�Kࠟ�����`���,����$Vw��<��1��T_�f��t[�ݬq!�"c� $ī���:Y ���NV3Ԟ�1��ι��^Ř��-{٪��m����I �_��N�h����"،ⲭ�n�A0g��V�\;��i��BE��ܬ=�n��yT��5@L�b��g|�<\N��YzlI�S��!�h�)�Sz�R�� �Hg�aw�+�,��ޛp�+(��߽���b*��8��<�p)�pY���Д]9#���k�� �_�ά��ת���rCL�N���Z��CZ3�Y5��v�q��r}Z��3Rp�7H��F6�z|�<�u]�����Grf>�,l�	NUQ�`�xP�d~��S�V�!8���0U�n5��3BȤ�T�N_fu��o������l�~31N�5[�2�N�8�w�y]Qu��ML��D3Z������bBp|'q<��w��ڢ|���z�aL&R�� ʤt�0��v�<v�J
�p�� O�=��F�����v!a5q;hB���ڼ�I�T�E���e�0N)/ >���F��@��H�<���V�5�\:%ߕ��vʴ���ﺑVu�f"{s@hO.�'�fa2'lN"�dW@l+x�j*��{N�Z�/����l(�ٳ?s��[�3���D�XB��T����{F���"[����GY��{i�_O%*�%~�e-��03玡��D����t�zCZ0��ٻ�1��8�	K�I5�>i7�ҶP]U+���jx�rj���0�=�a7S�0�E(H�U�ѻ��~�������D�.��I��1s�L�#jӶ{��P/��L�wj����t�D�0,9�\1Ϧ�.49������oP��t��Η�|�Ň���+��.�T��!��τ�xQ��F����� sF���`;iAG۹�t��H��^�i�Sd?�s+�daA��'Z?ɻ��
���yqF���u|\����_�׬o4���+5��a)��rW�?{I�~̔E����Όl�a��Ϛ3�|9_E��aLWyg@}3`��i���7���T�X�R��!� }n����$�I<����m.��[=�|��l����[s�	q��Q���&��D�PD�!� ��,��q�us%�̽�sU��n�%��{�S˵��c�$��S�󱵓���lD��'l�`���L�^���~��~�ױmϲŸb����j��IgsT�����"<d�D{����S����E�$�l�qŭkRK�ܠ�������tu�EO�X	��Y0jnn��������?8�{g#SV�z�Ġ��U6d��ۮ y�=�wT�y~��0V��oP�WT3C��z�!3��4�Q�\N�o?�?0�z�����>F,�o0:�ذi�`��m�h��v��Ľ�� dt?�A�I��~��!P������,�v:�n�y4k_��24��������G&������*9-�g�
-�d�{�E)��3�/�D�ѹ�i.��[�_F�����P)<˱���+S2h8��#4���2m�+�����L���8�I.�4�P1�HZ�m>.��*�����8�	8f��M�ξjo�-)́)�^�'���DC��?��A�7��r��*�Ql6�9�8u����0�~Ӣ����:���_��L���y��͂�����3�Rm�H9��Q�@�V}���/1\	��d����H�L  e-J� �e:`��Q����-Cn6	�rB;���y6GZ�|Ĝ��	��0�A7f�>+k�."��]c�ZFcv��
J�?��1��̈́K�lF�I�a��5�:�?z8����>zP��� İ<yt���ػMi��lߘ�~�a�HK�rFY?�$�!G۱I������s�9�8L�����O 7�H��B��z�
�O�`Ɲ�
��Jθ����~�}�ȷ�f��G�������4@#���D�A��5v��[�IBu8�ez�Q�ﺻ
�H����N�����A݊\�l!����$Ƹ�'���k`BF��B V�g�t҈M�A������plY�O�Ǿaz6�y<�gﳪC]RH�oE�VX�϶�;x=��Ӣb��s�[��%�6��¹Oε�]�ށc�5�CL��uz�?���$��`���$��h�6��]_]%�ߋ�q�e.�{�ž�֕�-zd5ng���R!��T�*ձ��l���]�-;�Tfݕ3_�ۮ�Է���4_ř}��9\'�;#�05��Ҏ��6��v�]�;����z�����);��^S�»���p��իI�M��������Q�Ŧ��n�1�v���T['�9&ۛ�GJ�V�_��E����Ĕ�7 �K1w�ȭ�͋q���J�j*�ԝ�g�S����O�Q�j�U��a];�Xwݔ�e�o���^dho� �B*<���x[��"K�0u��cw�VQj�#���П�(�e���Gffax$Eg��@��XJ�X����ȴP���t�I@N�!s��F�Nm��1��8��.DT襄�N䔯��0�"6j|R���) �|0mV�6�@��{*�>:����Ґg�����
xt�M���b"n��k9g��Է,��4�(��	�����y�'~H�o����\o�\j�6v�W��ñ42����vI�0��߸�_Ҽ�^;u>���Ʉn�;_Ia>2ɚӜ���o��L�dc�����n��uA��}�b�����~.l@���?�#�n<��q�����{\�h8���>�\��v1��X|Xρ���o��XT��\E��چ~�m��1=��Z=�� P[3e��l���*|��g�c��<���{_E�;JȮŪ]>2viE�V;BP��ic,���A���� X"O�ߓ�Aћ#k�>�����3�UH`�s�{��N-GV��f�=�1�����NxB��m�R5F?��ģ.�lO'�����L�2?�V.�I�f	��78��8QL��^?����)����uCs���\�r�����һt�����P�����[��ڵ�5�Z��Pq1�?�t�P���^1ɚ�����s����b��QL1���(gwG�)���iJ��)nyyZ��d�SK�l,�Q��Ϣ$b���WnR������pL$r��i�#�c`�E�����C�u��C�=��}�B�9�_X�<�#h��N��]�����5G9�)'�".쏬@��8�2�.t[ڳOհ�!n�E�.'�gc5�0���b�&+'��g�9=x]������U'm`Ԝc���s�ye�6�gJ5�*�0�kJ����&ֿ�j"�\���l i��>Nǟb^�Sd�Z��V,����~���ع�$�!i�s�2��ʐN��{u��5M����������@ꄫ@����4.�A�EN�� �"������MzǺ%��2G��E�}÷�r)b�O�YP|���K�Sԇ�G�%Or2�1�;���� ^3�T5�^)Z�U���v�������-7S�ؘԭ��q~�,|�Sp�Fj�:�
Զ8o?�O!�/E������T	��[��:��^=�7��,��8�����,O�L�Fi�-�Z��I3Q�N�r����`R<AR���Ѷ�\���h������p�/D����c��5�O�V+D��,2|&�&��&��f}���$z���)�7{�������|�O_�|���&����.��2{t#U��Ghb�cuR	*�����\�ϰ����[z��t#�;��rܴ֘ID�bo��&�{ڥ]���|c�TԠ��������pM����Iƈ��3H�22�ͭ�����|��MP{.�L0&|)�"[6�V"Q
�j��;5�����\����y�0[[��8����C�Y[�Q.E̙�O��ܥ����m0'���W�'/U�R��J�C#,t����X�u�	CJCH(���6X�ed��p����Ȓ���`7�5 1�Y`��i���Z�T��X�ѦS��:R���	���+�o!��e8�>y$ 7,���`���!\�Q-�LZ�kQ�\��3ݫ;�9���rߦש�`-v%ǺI�e>L�h0�EI�qqn}���y�*���]��pdg%bu:t� �y��0���R��QeY������8�����R1�WQ�9KG�BӁ�Gȵf~{��c]+����,8�*�"3}�Y�.^�u�`��7���A�^�ɞS��R�"1ር�\<�/�~5[t8��28|b;G�ׁŖ�0�M��(go�$�R{[�L�m�4���a�C}���-�l�3�1�%�V� �s�-��x�U�ƥߦ���J�~�3_�鴢�@���6u��o9>R����5f9�}[��C��]>��/�&�׭�Il���`ܭWÊ�f:\:���3s��M���_�h,l�lk�zU���c��r(蛆V��̅ yf<�Ӻߧڲ���r[kx�;�i�'<���~׹X�qw��M��Q�+�u�"~����g���%4K�e�Ƙ?Gs�W柊Bg�`��yk�G}��&EsR�U���WeH�8d�I�md3��%�2�`\[͕<Z��Gt��m���r9����N�A�C
���Q)U5�c��r.i��"�BX�����p�@����C
��%�;	�)���mv�Q>��;�:RO�R4��Y9ZW&�	���B�ЂC���u���ӏ��\�4��������γ��#�wN�$)P��T� �p��@.��3�4}n 1_S��0��0���E@�x�e,
��>�.���-��Da<�8=��M$D&�ϣd�'�zk�ȝ��+2�����:��I�N<�n/W�Z�M�\����=�<;���䕛�\{��X���\�#����-w��S�[H˔i��,����6\�y�n)AT�m]��H5�T܈筠��V�W:�]���^ �l\���ݨ����8"��31�2�j���[U���-y�Ⱦ�F�HQ�D.��!�

�g����+86V���8�ˀ��8�g��,/��b�	����3T^�k����t�.�AYH#U?y��+�eW�\u.��\}�ݺ�M`of	5v��	�Q@�r�W��ٜަ;&�S0k�O��Z�s]�2 d�tn>3��!�љq8�L:0����&��0�Z嬮��Sw2�6�ʜ�NdCF��v�X)�Ue�RGk��D�s (���!�R�0}ü+�t��+̘���;/�������7�)�i���Z��0�d7>"��f��J% k ��^ɭgH�0<�!������P1�\��5���t���!&
�����z�@F�7Z�[��5_��侣@Iw��EQE����IL��^̙���P2o?P����'k\$��U�	���k��߷`�r�J�8{����YS�sy(�WfHBmx���:�����X�L�h��ĺ�T�ׯ�iX=)w��{ �c�(Y>N�+��|ܿA<iJ�Ux�Kʩ��~��#J>��₥Tt�al�������{Ճ���GX�(&�� �f�����]󜮛�8�L:^xU�_Z��-e�-��!č��`Dg��`����y�2}����>�k̣�m3��}�uۥ�%$��g=�v�:r�T�U�#>dzt�2��֖iw����ߡi�$*�l�T�@~�lF8w���߻R ?[��yZ~��$9��j���]wF�?����#v���I��-l||ߌ�N��Tx^��8i>Z6sn��U)ݜ����)������D�m:�ǝ�9	-`�G$]�W^]�.;3�\т��9t����G��������9&�}i�nRi�E�R"%�kpk��Hy���h:ט�`�[A։+�ժ:N���@Nkq"�u�˫B��A�'�F��
�k*+zm�{��I~ͽ*d�m`�}7@�PL�(��J{?�a�Յa��-��ל�_�q�c������;Nx�	6�c��/L���\ (yq�WOɄqdH�k	fϵ̣�$��F��>)�";�����F�l$�й��Z��F�N7�������dFH�:`��f����G�zp����=b��4���ȚO��ế&R������<�tF90�;d���Q��B�����w72�]P�=�Cqᾄs�;��a�@�b��<�c���uh$x�Ы�|d7�*�R�Q?��oH�w���=�yʭĦр�2�^�w�qː�)m�C������?��9��#�d�*�.�2N�qǍ�������k���x{)2���Ç���z=�P�{K���QC�4S�0^�e5C*w�z"�h�� �Xf���xǚ`��	Z��x:H�Y�/��U�	��D���
�3ՒQ���?� MA�}��"i	�1�]������CA!)���8�F:iuF�����֊l�M��+}�6�ڹ�Tc���kA�$v9��hd�M���^�0�K2s�L����2&�+S,[n��f���D�\X��b�%g�6��%�b�O��s��{�f*n"���vc�}�uⱆ�a��P�A�p�.yE����:��R^�&�>�Ս�0ī�ZA�и��!���Aթ��������(�����X�̖ueOtSy$��l�����E���c¡v�Oô����N:؄?:�#d3�Qbal���Ҏ`X�����eʸac�a-�AF�HX]���ک�Xx�rh���~8�8)ܝ��.�RPs�*#�'��|B�NQy4���r?�,A=��wS�c�?x,�s��"�44C�ȎoDq�Y���W6F?�p�%� a��p���귗�;Pgkq����զ�C�C*�]:h_��2��	� X��+�Xܐ�8g��u����k5vG}ο
24��U	�>��<��|���L���ǜ�Ffjcqa՟F1��f��p����]�l�o" f���*�Ĝ�:s�Z�@�՝����T�^�`�_�& g��>�T��hT���'�YbQ��$]�Uk�b�P�;�u��}@��|m�+[�I3t�.d؆C
fNR$�5iz�Rv��/К�T��J��B����OC�9#�ڥ��3��}��+֠�쫖=�KA������4�����tll�p���ZL��)ɢ����ޠ��fL��	1�v�&�B� ٜ3�᧊�!����m;�eS@'Ř��7����u��A���h��[S)�K�)��3pׅ,�ů[C�#Վ�8l�XlxVHYEB    fa00    10c0{Uc��s4����7m�H!�THU�u[�B{D�~�Fb���ZC,�Q�LN�m_��˒�Z�����\�!O�˵�n� ����ߏ���
�g���Ns0��Ҵ���b��c(A�lJLk�ֿ�zWl/x.&@�/��4�Df�m�뭕!a�8�#YGr��DQ#͉G3����i�)��h��R/���q;J(wf_M;��c�5{�aO��bZ�������ώ���G0M.9���iQ|�d�|_p���_�N���v���D�9Pc���Ö����0Q�����M�.�u@yQk���ϧ�;XT�+��@k�0�b�@�������ԑk�-�!�l/mK���k��mWJ*��H��!�_�4���7��Ϯ�e��2х!��9��L�G�SџqP��շ������B �7{����::���Z��z�d44�&V�A1��zWj.G<��/�a�;9�>�3�$�FyRi��HO��)H�VE;� ���AY�G/-QF���Z�+�w�q�^ݻࢦ��[�����9�C�|��?�%��S�������$�����Ͼt�W�E,�C�Tz^�ߞX	τΙ7��µ�ql�m������̳$U��p�^I[9�"-+׷=x<I���ȑiv,�}?}[����b,��È#w�����,9����
R0�����ҏzُO$:��t�����Q\/��QUoA�-�h�"���f��$x��\=�뉉�T�}��߶�7~ط�O��x����Ih`I���l;%ȤVY�Mj�<�~�|�Y`t����QQ�/�ǶM�h����ӎ�>uH�d��_1 8���&5����~�%���^z���;�=�,%�4)	H{i�p~����r�	"�º�5\;�Kx��l�a�CS���2�|��;�5*�%=�3�R�o�Q�:c�0H�0B���w�5�R#��i�﹚�.�$�Q��0z���c�9���Q�I.��g��-��>�U���yK�����x5<�\G��As�L{�� �$QxҨ`jn�$���o��.Y����_;<�\"�-��fݕ�r�-~O<ڤK��!��^N���\��{���O^&4"/�/E��S����z���v�9u�c��������`'�{m3R��kg��f]���y�p�BQ���&b��v�@��i��Aw�����-@N����zSk�}�}�'+���U�[3ɶ��9u���d� 7��������X�wT�q�kiu)��>�L~A^"8;���M�~2��-�c2�cQ^{���=�90�����=[�#���T\��u�LEi����q��ꠚH����x|z��mR��
�{R�T�z�/�B�쌏���|��m-?����A�\�BQ���Z|�U��x���r�/Q�����`����o�]j3n��w�XHp�Gx�vF�9FZX����G�1��L�O��=��p?����.�(���������cnџ��� C�R�<��OKE~�E����>��tM���+M�ٸ������h��:��NK ���F<5�_G�ct=�a�����}y��
{�����R�oŠw�O3�yxD|������7"��^;��Y���ҫ~��B&�x�ΥI�Q"�cuأ+��zɪ�="����!�J�2��Z	����5?"�_��ֳ�Űv+p�����l�`���S��r�	���X�'�,EH
΅�XX	r3%;���*{��ݭ\��	&��u�;xu`*���_��Cs��2���*x$4-H׃�U�c�U:�& Fb �Zi�٪�u4l5c.���s���M;��8�`�@F�txBQ��c�UÖ�٫f$�;WF&&\W4�(�챪�]1؆��@���.�6f$c20�w���<H~�ZT����O�	y�9� ��&�����w���vQ�}�a��zi_�������/�x
��q�C�+Ԙ����8��oL1B�%�am�T��N\Lf6o�z�"$���V�Y6�c��:�L�r��;���g3���A��$ح-�6,�����]�]����y����.�_ۀ�	��9F/T�_��/�wz�_��̑և��<2��+����&��.�,+��' .TSsL���p#iT��+���]�e�.�@�J?���dnӼ܁F*iH�'��v�b^�ʏ��8Gɑ�,q<B�~'�o���G�_r�L�-�`��u*�a�b����Ma�S|�s[;+�0>�e�p��p�O�=�nt�����;��?��W_��W��+�P��8Y'��ո9O��c� X!n'[n,�y>=��Ҳ
~Ö��Ns`��V).	��b9R~����v���Pݨ|\�@�����G��K������jKmn\�؅>�>B
<��צ��Tj�L���AyN�\'�qE��I��"�� �O�۪(��6!C1�����*��6�5Y�7^?m������!(�
�"���]}�7��]#G�r�"�l��`/��I� /��M�&����TV�!��$���*Ω�-�z!}�:~-G~�£ήr��{S$��G?5���I$W���[2b"�����0,$?ŀW#��Qܨ�\�:��ZY�~�#*�J�@/M�����Ig��J�$��+�[ 4�cՀVJ�B���bm����	��r_j��@���QOX��-���$�� 빉\�e���m��]#��py�T�"�jd�wA�LMσO��g$0p{��`�P��l; �aNJ� +M)7xh�> -7�Sh0�����L��jQ�R$@s%��Stl1��`�����gYM �|���@�d� dS��Q�*�ǆ:5!�32N�Y��=��bL�'���������;�Ih��:O7XI���]����כ�z�;�{���[���;�Q�OJ��G�;l@��}R_u�V`�V	D�Q%����aҍ���~�1\�ϩg׆Tc��W)���/$�}[��3[)8�܁
�&�?|N��dfcB6R1u�6]�� ���ȣ�D;����1��1�@�%Ƶ�f::�,Gs���?3�*H=�R�Ql�xgP�gHy*�y�<e�9���-�O5)��5\��m��麤G'�f�@a�-�)V<���|��C*�L����3��ʧ�d��kRq�UA%�L8��!�|�x��+�ɑ9�&������8u���hɱZ�����vn�8��ޝJH�fc��gx���"2��[0h_�NjF�E?O0PQb�����m %�vM��m���������K���ơ��n�n���O�:6n�(u0�J�I�c��&��sE�hIҩ���5z����&�)��I�r��,|�r��UK��+HX��+�M���u��H:He��>;�H'1��Y�jI�����b%a�Ɇ�����a&q�.}]��rP��+L�hŝȻW�gX/�ݴ��J>p�'�\��o��bӡ�@���o��m����������0���&p�VWP��`KjP;a����F�f�C�J��� ����_��9XHO�m���D�Q������ȅ���W ���@ǅv�D++ޤ^oQ�_+�E:ϒx֍��7��Jz��/��dn[�覹�0�����{����N��U ���#�*z��Z$wk-����)��4�FQe��A`�%-nP�~���N���˵"��&�kӅޘ{^ Ƞ��XkG6���9r���:�K䭌t���4H�^�c�0y�~r5����*x|���W�A!Wٻ�Ń��rQZM�E.�*��U~X�^n65�^g�ug�Af��� ���&� h&�P��5�q��Usb�Z�-�[c�?-�&6̍nO΄��5?�7G�'������QraI�����aH�-��� � v�ج�H]v���&���0M��y\j�?���+������趄'VR	Mį�ݗ�
�3�{���r(�1ʴ�#wH.r�}�F����f�~�HL�T�� @^M���M�[N�K�XStP; ���8� ���-�.��6�KUq�"�\^�~���D�X��߭iJ[���1Y��X͞�̃����oc��κ��xho�$�B笄��	����� �&�����K�}9vP��]�c2_R�@q�0i��͊������(�jHsEns�A����|.����z�U�vh-�O�(���[?��L���{��a��Ĭ�3��bЛi���=��8�A=_�x*zVdD-�|З/#�L��	��d�J �i��D� �J�XlxVHYEB    fa00    1140��	�)X�jo��~��X��R��x��t�(Fx����4��U�B�&dk�p�ۏ�t?���S�2`o ����Q1F�,�(����f�ޛg���(�ϟ��������%����]�\���~l��&p/�5��a4T͹�H�%�ě1u;��-�e��m+���n�������^U0�}�G߫7Kצ�mL�	��s��y�2���7}�]����h�a�գ�|��ؓ�ǅd�)=�n۱�_�.j��x�I�[Bl��!ba��,�i.sx��!�����7�2�N�̦��T��8����1-��oRW�'"�ޓd�ō�<}�^J@cT��?a ���_����i캢�~�$&�b�z���$����K	�dxX�>p;��̘�'��-̃"����67�ˠ��RLw��vrQUr�u俷�%���V��S�=�:^�7?�|zݏr�3 ���/���Oq�����1�,ᘓ�H����#&B����pRPӶ�M�䦫f)< \'��PhW=�{��x(�.���ԅKǚ�E�9oy� �o��(��J�� ?4'�.
�C#iH�צqlK���'k7À��v�d��Bjog�k~��9�Z�Dku��A1���@�F��P�~�����ݎ%���e|p�KJW�fǑ)��i�.��mǣ",��ٱpQ�n��|�'�*a���>'�,/�����=!i�0�hw֖��!���ε�9�H4	�k��+���6��Q�>h;��rd�����زŢm�4B�э�
=u�!�t�m�5���QI�n��Dw�����P���T��x�1.��B����^3����dc.�V���4�r��L;͔D��'˫���V|��S�y�B&�O�-黿uy�����Йِ�S)�_%�x\�e["��[|1@bz���Y�r�EKY��$]�l����»�و$�#n�/�Ӎ��S��IB[S� ��H��~,@�,�d9�l�S�Y��``��� ���v��n6�#��^�tJa?�`��e�����gE�Y�����Z�%D�M��0HzZ?��ף�~�!��I��*&��h-��A�˙��h�Ѽ���(�Ȗ�Y_��η	��?<p�GD��q0��:�� k
��n�UQZ�X������
"�K�$�D�sB������ �C�=yޥ�`����/�~M����^�,���M�ֆd�H��:8ͮ�Ob1�:��~��Ʀ�V��(PC�MO�"���kz����}R�7�}gx���b-~�@�+����K�bӎ�mE �?�����$+�Z)􁂴
u-�ǄŽ�@�UM�7e^]�:�Q��G?>�Y�i7�P�]"G�n�e��� *����&5A�<��@�Zs�]*�(�
��e����uK��;,�=i�|��$��b�����C���@�߳| �Bv���M(=K:uWE̬�S�q	�T�Wlǧ#����O��\��2'�Y�X�GO��f�=�)A��]j���S�F�wN�ˉ��}(�w�&��ڨ�r$�'.�Z��@���0��-~3�d	��C�D���������p8�_�z�1��s�l���$�v�eY{|qt#ĵڼ�ێ�L��@\��i} ����;�b̬~��0�]�ҡ�=W�R�祬���R��_��PK����:��[*:!���X���Ԅx��{]����PF=hS< tR�u.�ʖ�
޽�������@Lr\��@��/�_�����A~y�����֮��(�(�	̲ngͲEj�l��i��׏a�)��EZ��w�|�@%tve�[�������ܸ��"��A��˹*�\�KaW�Sk���I{p煹�͞�5�I��.�A�C��H\����e�,n�;wp�xQ���Rܳ�L����0U(jW�V5��τ�UM�����6��z$f�w�x��<
�.���o��������H��=��8���3TB��f��!!������luy3Hw��V_��7�\d
��v���q#v�W�]N�� tC���V��H��R=/y$�"��f�hR'����W����g�f�i�G��5�6`��F�򴘚��0�� �3,Ț� ����kG���MDz�)�c�Tō��-p�jإ��ឥ��1�|��{X��k�3�g	oJ4�:��B�3���a̳�J=����U�̟���	:M��R����ډC�>��a�Q�l�d�f|8�D䲛��z��$�;Ѵ����o]� ���z)0����il]0�	�� I��{�R����.�N��2�Z��y�M�jw�?�{��{!.��1�t)~���d������'�Z���{�l[#d[,�g�qNAt����́+6~a����h�&Na�C�����m�m�WgW��ƀ���I���~l�%?��<yν.�����U��J�o�3����O@�CB#VWr���T�϶ە@~��� ��Qx��*!�g� .�a}���tf'$�.ǳ���%�P	���L;$<5i7�Փ�e�f�H�8���B��8�27R]b����+�A�Q��Ȧ��*̗E��+ZT�K�,k�HE���u�Bn(�h�j��9������2�o��h��Fi��k=oR�5ESM@Q
΀�`]9�wYY�
�H�v��9���)����K昦���o/�C�K���i�Mc n�DIzN��"�����?���W���]l� �i�m�g�<NZ%�?nb)5���u?��o�q_tS<4�uCD�_�S2����7�V8�A8�o�������X��J�m6n'�(@�|�7��җިR^/Z9|W���GI
JD�2�
o-z��9�WQ�U��<��r�#o M�m�>+'uȁQ����s��1���aII-?$���C�_N�Yw��V��%�H�0��3���!�4Dkf��˫��Rl*tAJإa��:,�}���[����C-M�H s�-i5ED�l�M�u ��Y�B����[3��"/4ru���<B�K1�X1h��N�k��5����b��e�Y6}EM�D΢�X�	О.Zy:�-��ĀA|I��BJ�1�>D�O�i����F2m����m<Ҙ���ܞ�?�����C8���R�����T/Es�!w�U��ԭ'D����ј Y4e��Oa�]�Y� ���w�� ��N�L_�7J�zQ�����I��&{�1���bƍ���-��y�{۲�rq�tW��R�Fx��/d�p*���	�\�;�!�P��\=�w�\E���"��=�����c=�tA����T`Ay�}��:�%���'�X
��EA��ڨ5�|�� �{�-�r�z�}��U]��������J�y��5-l�_xKI�t�)�(ә����{7�]��rp�W��Fm����1�d��w>Oν�YIZ�w�������٫"Xno�����gJtϬ�]��JR�������qVr�I �����F 1^g�΂Y�k	��?dhcqM�Jk�$|P��b	�Z+��d+�@�x;̻#z��ǤN#��/^�ȲG�Z��0:9̩o�=_q!R-2tm�qls��]V����%�/�p����٬�l{]�ԇ f���0*4yN�v�ݽ�%gS����_&HC����]�	c��;U��3KC@7��\?�%e�,���z6��΀�_��X����y2��9�~go@k�ߍ�|�d)�����8��RȞE��j��^_C��J��}5,��8V�/T�u	2|��9~��ϑ�D��_���f�8��ʭ澘域#!V�ܤ[�G��Pj���'���tX���yd���|���$:|O����G@A>�=i����v4��S�����|H�O%-X��n��5��w�ci��7�rc푋�*��{&m�ptD"������ٛ9���sV�\�H��6��'h�x����J-��P`/Y��Ϝ2�Ab�e-ty�Ҵ���=��!K]���ʪ䷝~��٘��r,�N%O�.4~2E^���|���}�_���6���Ĳ�\(w����m*ə�d�dt4�T�ݐ��O��E�F�c�����એ�
):��"U
��hv ��5� ��^�F�jB�H�:%�N٤@cY�!q<��:��d�
��*���C�O�&�K�/n�;�d�@9�yoD��@fQ����%׆a굛L�6)�'pAM�YQ�N���a�E" �[��O�΅�Tg�я���n�P���|�!N����۱{�OA�C/�7�q�Su��C���"5�֛�䨎��E���=;8?R���JH���%UAK��ؠ]���<pVj�$:=���(�A=qgujXlxVHYEB    fa00    12e0!������6��V m����5ޢ��N�G�6�!�L��9�T��y?�͏���ahA�;R�{���#�n��Dc���X���b��d߇Xʊ0F��0�E#�$�3�^����isY��ǲdo�f~�'�֢�^�D&���hu�������ȳ�˔xg3?�q.�)�{J�1	i�)�����-Oi��p��b��`�cʓ��y��=>]E��_����\�T�tB���4���8�oIw�S�9���~,�9r�d�̽0<�)R�(o�J#�6J.����{�����ܗJ���ޑ��nط�=�?���pNM����s�c��.����k�_�����l�3���-1?�Xv������U������]�@\���E�?���~p{n*(괠z,������cDx��8W��*/P�PoXL'����|hZ&��fF*�mi��oOfi^5&�����qwdz:����:��)�.�~5��0�PD+V͚{H�!@C�PbN���J>�H�s*���W�	7�RبM���}�$��9�=��� `�m��â�J�瞩p��.�醤�k���k,�	�t6�_�#N� �e�6IQ�����6H|5����h����:[�A]���Z|5s�j�<ϫ��J .Ȗ��3������ t)~X��MD��bG�2���Ԟ?;�)Z�ԓ���~ף�6^_����<��@��bK�r֟����~o?�����V�M̈́>N8P\a��@,H,�l�^ ��p�-�Պ+f�|��z���1���5���\���?��'&�bM�O���gI;�V&��
K�{�aTˋ�4��|��1�"�ܪ{2���&<���ǈ�_�uCE6��|�����+EB�EZn�[���\gn0��� iÆ���{#�%o���@~��/��&��h�`? �]�C2��!}���bOe��i�AG��S��L2od�w�k5�����AL���ٖ��hD��>H�h��E`B��g#��;�f-M��7����\K��ǌ�&9��������2���l�z��W/H+5� 5��ǆԸԈ���#�޶>ZUM�|TG1@���<R?H(,`����TV
�d��@ez	Է�~b���\�\*,T���5�k��0�� �H�q
m��������p���8�;���ϐ��oq�1�b��tX��W^���oF7��K4�����R��� (d��rʉ���:�;��rE_�`?\��Gg�����8S%�,,+(��G6�B����f��}�����HH�zEFx�-*�����(�!�l�EޭL�M�8Qc.�{-��e�S�Ht?�R+�zQ|�&Q1��(&�!'�ᲳU!�c�&�а��3}
C�ɿثF�B��+�M3]��/���-4�۟�mV��|��)p��Z͊ob��j�T����nM�OJ�����o�A��!�'Bԁ(�0�<]�'~���&+g�� k�i�c��eT@P�y���!,��'�����w�!8%V��hY;1{���a�Re�r���8�.��3�15������)�5[;>tؚ�ۄ��;Z��t���ѿo����*䓗������ �(Z7������S��S����/ؐ�)�3p�
A8`�C=YOC(��Ŝ��+�o�w�z�W�@�,g����ш\HP��}w~���] ��~0�r�O��,�j��I8��Knqc�*F<���'�����d���G�D&C�pb�Q�rr�gM�hQ5	��bw�?��"Mt�-�-Ǿ�㸝������h�.y��8J��q
���6������3�����x��"���)��&�"����8ׄ6g� ���Y�wz�g�j�Ɍ����}*����0����~����xg��
��F�ABq��0��md����$v1m:HCH\��*
7,ѯ~������b�K��4_��b�h1�072���cN�)"�]�܀��;��"���|�!�:��%VO��?]���̏?��ސ^J�R|�zO�|��jȑ"�7�7sQί5��pM������7��R�g�Y�?g�_H�Y��x_`*e��n��y���&��Y;̑~M�Tl�'�/ڪ��Vs�߹�=ȭ2->gU�v�2W:����W�6`�=�j[臱�0aLQ5@Ǭ7U�8Ą�:�Q����3vXLL̻��f'o�%�D�8.�}+ۢف���#H�o���S^�o`	��oI�=fq0<���eN3�}���O�w�^'�����i��GO��� pm5����'~(����T䥘{��b�AAn�p'�XA�$d�[�ӗ���N4��B���̍�e�}���<��G���er=b��_��`��c(-'�1D��lle��-ǋ93{I;r����������2d�I��l5Q��v!�&C���<��nV��>�m�2ë0�@�Mm�R���y�w�!6f�JPI5F�1�0j�������eC����.Y��v
?�?�EH�0/�sg��#6�	kjHtey^�@��(V�\��-���/G��|�U����Ɏ���X5~Vf/�:��OU�ĵ�M�S��L�o�#b����$f~f��.JK��꜋k	P?z��x��f�72��@�p/@Y\N!T��O9t��̓����6�^��x��u7�"�<�<�^�(ÚUռG廥D֖n�d���/�:ǦY��b����>��gsH��Z�x��5��'	J*̽�� ���_�a�|�O�%f�]aB<���'�53k����^[�XQ|s���o�cc�<���r�pz�*���?>��=4��e��J��l��m���c�q|�IM���L�O�	�B7�������`������禾��'�X6�y��f-��k�}-'��*}���Å�����|\T��a��UW4YGɏŠ%���|g܌��r�$$�i����ab�Mp�yf*W��Y�b�Q���aϕ��!�)�s)z�m�s���Y��A�"��R��;�8�tҶh�,n�˩��߂l'�tt�t��g��cK�O�.ݑR��La��<�=o��e��BݦM"LGDc�4%�[�8����*u�yF@7'mٖ�Z��>�mkCcgK[hD�9f���j��T�~�ph �#xka�{����>ofN�?����sC=h5^�T��Mg�k��Cc]H��Ao��\x�q�S����Y�,���V��H��~�?ƀ^>]O�b%\�8V�bȠ�D|~j�����?�p�����J;�A�;�׮����zy����0�ٓ��&{��̲Xpg+^�tZq�"��V!��fk<	�6+S�P����b�����w�{?��׵�����"]'/��������to�W�PkR���8PN�T�i�gٽX��1�Ix0"��m���o�<`"O���"����`�;�1��Ő'�/�t�f��ԣueoF�@@Way5|���x�O؊��AM!�Ul�LM�=5�v0���N��Uh��8����KA-�n�"��Z�����{Riu;v����N��y��2��V�s�@�A��|���Y���JR��ŵ�pK����\B����jni_��Ő��t����m*��p��t�爉��.�OU��5VJ�+Z2t
&9���$���1�!�_f�jS��I}��Tu�.>w��y��z/�N�\���V��~h	��_V�C�r'�0���{�)�ƃ~�l�D�9�x�����h�ײD�m���g�������8�!�nʩ���V��X:h
��A�����t�[�U�\��ƅ�USȒ3�v�I�2���L���ձ
�jL㘘��҃~'b�@�Tb�d�\\pA�4p����e�ڹ�#.-^���ɰ���LW'�#�j��O�k=�����
�C�����F��"�[ or'j��H��Q��	:��kd7NEp{ʍ�%l=|A%\�l\��Kε�[,�����T��s��u���v�?5�;a1����@*r�������#�����ϳ��3�_��rw(���,��ٟõ���C&�k��,<-C�b�_��?�YK���&��e��n1���'�څ�Y:��0J<]U�j��{�M�PR~�0y�gKw������R�N9���E�A��V'U����+����Z�a�?=�w����6�f|@9���maMMa��H{���吆�V���/@��jk�~��èV�A���=��~���	��XԨ8s�cqㄭ�?�9�:�}�����e�gZ���2gV^�hE�J�Y�C�\԰���ua�#=�(�����t�Qx�GK��?�*l��j�=6���o�2\P%�-��6&����
#%�Y�����0)-����7�ن?����1�8�ҥ}=Wڱ��o�g�i�7�AхP@�Q����`QqՄc�⻣��<�j7dý��?����@~��ODP'9Ra&��"��B�u���=�j�3�z7�r��[�"���]|s��j��r*�a*���z7�;��Q�_�..�Iz����`�;��m��[�E%�;X���{��F���^�LkU���P��b2��8f\'�R��4B�Ңbb�Q�L �W�������@':P�O���gG��Ǒ�sުP���o�'.{&�~�����	��|����e]�_�:��ʆH�R���U����r���9���P�dӵa��1�*w������k~��������������ͼ�D�;�Ox���*��g\����XlxVHYEB    fa00     f50�@+��#�~�7nIg�W"�����9� Γg:�6���1��4�f��:����$�+aeAk��-��D�S����I�4�M'�b�"gA$��n?��G�*�@�?��I���B�
J��!-�<s9v(S[���"�l����=b:��h���4�L`�Z�^	�y�;蓿f ���庲�ן%eJ��v�8�JA�����;H���P^��yQ%�9��fS���r�u��-��5*K�Wyac����SO>�Ae_X��~�훻�,~\��˘�yfB�z�]��8��9G�#���I���Aȧ�˴n�s��V ��G-CF8�%�����c�
� ��_Z�<
�C�z��Z�)��)��V�V�Q폒�j�Z�U%A�v���w�`G����0N.m$���N�H`+$�l(%
�a��2�.=z�u�%��H� )�{������&g���E}���"��S�+N���е�w3:Ь��~��sݟL�R�k�(^UKv�>z�\J�y�$�2��uS/���je��y���3M�����~U��=w�z3���k��ͤN�q�Yg�$�^��׈�!��o��wؓA���A�-4���z�xe�[����:R<]g��p�t�Z���X���x���>>-=iٖ�xI����	�Y`R��w�%߭�m �n�Bn�~��ϔB<�j����T�ZM�5�	|�L�B�QrZ'�F:�DX�fQ��.Y��ܦ��������,5�DzᏚ.g�]HM{l�;B[��X`�^g<v�F��f��SQ�������M�>l��Ό��I�)A4ʍ?u��R�8�?��[�T@�kXhP��������Q~��LCK��<Y+��rn��0�pK�g�u�*8M�>���>�~*�ܫ;�����/�]�P@,F�m��r��Q��_B]�Ś�d-짷��w��v�zM���-�D��\�I��#�t�~�9��4�<d��:1R�Fs�7�����<�"?ѿ�jh�b@d�Lx6.����6�[���V�sX�-�m��+�7|�;�bSyUƸ?2�:��T�#���p�2;FE��k�=�!��0�#@-�2��OO�شl�|@��f;.�O��/���^�9���xg��꩷N�����+���ش2O���n�S�\bi���b����[*�h�3i��DJ�\^�=���XP�k�O%��'��G�~�"'�A�6P��[���!���|�-\���YLs�������o������l�{>�R����9?3��A1W#<9��'X2���]V}������*����z8��
d�n���#�v#�2`'��ϕ4+��U��ƋA:�Y��_��BZVJI� .�zu����#�II����"�2Z���B
�! ��|��/�� Zv��slӑ��TT�5�dU� D49)�HK����,��e=��p��+b��H)��j���b�/�$�'���t[7Gi�Dv,���� 8at�"�Pkoc�4t�����/�h[�ײ�y�Gf��j,�^E�]ʩU��M�F!��"�2r?�F���E]�Y�3��dI�i�xa�9�j�K��&���)Q�΍���,t��1��~�|����Z�F@ƥM�p𢶆�F�ƾ��A3eTIx�➅�S�;n��I�'�Μ6� ����z2��3�5a�86>T����Ļ?ϖ��NeI�0ٸ9	e�sΊ�o�!�"��'��Ls9-��Id)�i∛����VC����t�y?z@��6p�5	GQ���zu�A�3j6�I67�ՠ���Z��;\B�.P���XV�	�s���^��
��b�m�d�G+��-tm1�Ƹ?A����z� ��=|��,��>�ZA��_��R{쉨�u0���Y�H�+�S:�S�w�؋3����|A}<�<���l�$9�%!Ev٭TU�& a��=�wmZÞ��UAK ��AeJ��W���1�w�}���#�Hb�y(9�p&9Je�d9Q�Z���y�J@Е�J ڗ�G�Іu��}h��Ğ�j�	X�;kx�*�?4���P!�V�	�+K5#�*N�▯���`@x�:���j��W��>��N����`9
\��{�6�b�K5J�a^� o��wv�ȓ��v*���o�0�ƳvdHid��:����o�������d��9����R2͘8;��Q���DFD��汹S�9ֳn5�p�����8�L�{!7o��E�@c����Ͼ]�&f�y�I�Z&������
�%3p�ے�z�J�[�j/o;?�s���ֈ�HB�[��s��~�<u�5���t���o�����A�zOhFwP�Riگ1+��D�,�T�.j?�	4���e)fk�D�G�q�y��^k�'��Nsho.�b�P�7�V���]�'��z�?~mjG�l�U��:�R^�J�2�(����T� ��ס;*�I��j)����NZ�Ӕg��K�j�ã���X�
F,�o��X
1'u��e���xВ������&��؄�����W:��j��V�.�(Ut��������i�!��s�[k-�;��|�Y���Q{��?xn���i�0~�WCV=*�4�F��)�鳴��'� ����I�^����g@RY�m�G�f���ey��^G-�p���0S�aË�$������L8�oBS��6�H�rR ��z���aE$����B���� �*�Zl���Mcl�HF����um�5!�}|��*��SH�
{�޹x�6��JN@���e��sJLG� ?�ސw'��d��]�N�>+d-�~ʄ�o�о�_�*0;��P%�uߴ�^m
�%r�u$�v ̆�{-�o�K�y-�
H�E�p�%����V��cS0�s����/���&�=p�o̗�@ەL�$��;%���q���S]��1�_�B���+S����|���-x�I�^ o��OjX��4�DD�a�l8K/Ԫ}����*�ܧ�}t�+�N������ȩkS���������O��o�./7�ߥW��w��%E�u��:����$�#g�}����/� w��I��^2j";r������I����7ҍBЍ���9e���:莒;]�/jyE����%����-�q�NO4�4ɮ&.��+L������u�S|	d��G����e�[�y8/���:������.�\��W���a�'�+č��|}�m82�m�~�>A�pUx���&�?��N�>��G+�x�"������^M�=��K���%�@r+�wo�k�2��{3��R��:�]C�*ʹ��ϰU��\WV���������F���Qk�m�\yz��e��+t�EF��U춠��_T�D��l��]�r�+�C��)E�>��*-�3�����rQ���ou�����qԋi�f�%.�.���,s*�"~y�d�Aӝ�Lf��%O{�vMi�ןR�^��AX��P0��7�d�W ��l�����x5*�p<r_Z2SW4���������>��J��C���z�4�LdTA\cC$H�(����L~��j��Q�:�ٴ��Y]%�,�B������5�}$l/_p���Pa�
VK��m�v:2�q�1e5�R&pFO�{�r��v�����t�`�s�/���y�S�s� )�4�)�kK�	b�*-'i��|��Y
g㪈��͜��L��w�|���49�2Y��C���Z�Ę�����b���i��I��✄i�o0������J.1y"Ĳ�XʺY4�y�Jt�
T/�f nNþ0���m0�涐�aT����+p���@��xu8�rP��	��7��i�g����:�oni�^A��{&9Ȉٛ��^�$	a
Rs	e3b��פQZ�	O�^L��XlxVHYEB    7273     560�[n�r8��ݰ���_�P��C1'�����yM~��w7�Zի����W"ms/9L�p�-_ �~�S�O�H�b��1�9ۗĂI|.�8n�l��)�+^q����]���Y���f��iF�& ,��AJ�P�Vm�~�<���ٸP'�a{f\!��|ϡ[�����3�/�S���2"qbԼ�[6�g���w�L�V�l9��+��A�����vYq�%�)8ْK��>2*������Dy!�h
�)��qD"��`��<ݑ{�#ᦋ&r�&�	�<+s���i	7
�w{���7ս7�%��]nP��oa ���φ�� �h��.�uG����h�z���#l��,����Kr<�{�L��ǐ��?KOAR�Ä3���\��d�H���q7+R4�n���y�+b��;���i	��:J^�o���{�I��B��\��>��}D�^a�W�uv8|�#��3�TLzP�}����r��l5���&���料5����.������$I�P\�e���a�����н���.`� W�_0iA�'��맶v�����Z��lw<��m��/q.B6���c�	x!�N�������#���S�^
��������}G�ݸ<���e��yo$L�8�^,{]/��W�F�gu��w��$���~� gu�Р�m%����T\ >ݢ����Ҹ�)�я��&-z(P��G:��YS��� �C8�h�ֹ�j�S�I�1�&.�������\��R�0U��*_��'���	�[�~=GLp��8�����L���Zqf�{=P����|e�|�:D~�T���^C�;��Wh��[��~]��(������j��l���0F�j� ]����t�j�*�t����o�`��3�~َo�=��=�����d�j�O9�܌���G��Gb��v���j���9���j>�)�˙������}�J`~�xK	�M�,��Œ$x@�T�|ֽ��u�B
H��}&q:�49�c�U>W�claW�*��+�,�DW
��+�h-Z�].C��g�J_@40��!^��?R �����Wn�����5�L��Q�gS�"�+�_k�<:0r� c�y&�D�w����p)�♼�h��)�V'D���<;�A�E�A+�W$��~�٥����4P4$�|hm�-�5���� ��<Ĭ7�x�5�~�]�s�;�A8~W��{�m`Q�t�QG%���`(@�Y���5Ra��?�S�/������JΫ��O;g�K4J���G�,�.���n���=_�2�u�ؽ"(�Mza��t�"LB�t��c;��!�d�A�|B�h�h��ĎJ�O����� ��B�����=⭇�@FU