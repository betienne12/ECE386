XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$���\��8�s�N`0Ae��;��D�}.�ҡ�r=�sU\�T2���o����M���#�W~'up_H6(���u҃�SN���,���w\s^�:�D	�D%a6t��
�:V��'�<k
T�oH����w�D8�]���d3�m�љ��kt�:�w }��fd���p��uLC[>�N��@8E�X�� �������A�)���ŋx�� �
�@���K80�"Rg}�~�e7���4ȼ���!�M{�춭$h���W��̿�~v�E��؞n��o��4*��YT��a�8g��vS����IeDP|�@?u���H?(��	c��A8D�����Oqz<@�@$C$�_�\rjsB�����b�Zh��{v~Q͢%K���3�J����y&.�lr�/q�8��](��	6yD�4�c�Y;#�?�Ķ� �86�9�ad�I�g���[��&0��?٘h��N����O�-(D�u�=���u�V��?�,�}d��!�����8C)���޾������*�3\����+��qI�ԙ%X
�м�E�|���RL�k���U�~�,���;�$���,�%o6.����>�}�߲�^� fQ��V�kh%����|ma#P��/��  l��U&o���9���?�r�|3���^冐`$o1+�b�6q���2�'���Z`���3��"
�[�O,s�n�Gw�y�Q)M���k��M,�DQ?�sY'߄E��!�k%�����
fS��XlxVHYEB    9732    14d0��ja^���/|x���=�x)�W�M�\�9��:���.}*_귴��k�zC۵�VF]�i0�*��BN���aCmb���/�Q���$�h���������u�b��JE��fa�뒽s��ӻJ�5T��?Q4A���91b:<o:�a�=y/l��Y��`�="�<�	���a�Y�%��-�ZS����{�� �+\	��h��V���'���O���킭;t��!
b��C)V�*�o�CqN?�N݆�'G0M8�fj��$�� ���b��ǎ��g��TL��e�zC�YA���b������.)����O;���uO߃�����]I���.J�Jqۑ˭զI]/5bĎ�
E01�(���P&�@McZ�I�9XW��dۼ	Y>� J��9���r�-�Ƞ� O��eA�(���z�n��Y�i�F	_#�C[� �RJ��H G9�����$	Z|?˓�b���\�щ��B't��j!d(7�ô�˟��B8�.��A�@UV�"�6/��m�VL��x����5�� �k�ϵ���5��D/�v:�#:ڢی҅�=$a��I2.�S����.8 �������1��v��>�?_bغs�������#�Q��p���WX=��7_J4�.���Y%S�b�8�5@j��3
����'�������k�F�U���q����K�"ȸI��4���l{�L�%���-��i�8�"�t��)����վ�~�� to���l?4��+@��Z������8|ଉ[A7����g�~���?���#w忯��t�f�:w��.a�Wx�I��mHԝ?K�\e����������֤�<�@��疿�Ͷ������J�c4żHO���� �ӓ*�����6�%)�����HF�@B�Z��j
j�j:�b���Q�|1�0-���7e���W������F4�$B�g�S.ІA�ܔJ�l K�bl"1��x݊�'�R�2�?��}M��YC��!@F��T�s��756�a������Ǔ:�g�].�{L�F}�竿�Ҩ�d��Ӛ�Y�~�c���͸�PBV \�dmbZs��Kr��8c�`�dl[���p�*uG�;�T�6-#Đc��va�W�-������ �A�����B��D�s�
�������J�rC��)�ذ��8�#���_��)Qj�$ �P���p#�o/�P̝z\�����90�x�}�WS��͏�]���;��6����2ٌ=�7Mrt��U��AB7��L}ȋ��B3��q��e|3r�
����%���c?*̿�+�0d�K�AgOE�BN|�� 2���%���E���لo�m�x��逕�$���G��G�e���X{��iz�4�/���
�����9�!96���nc �cH������H�?�6T�cz-��r�t����t����}�p��2�dޑ�!�_�s)�Y3�3�yp�ॾ5���HHݯ��3)�Њ�a�~�i�*�f;2��8�Y���y��<��D|&8�ٔ"	���H�X#�_�Y_�[I�"2�cy��\���&�i��PW0(���;��ѓ�ܪ_���#�x,W�G�6�D�&�΋�r��4�cʳXrU�\�0�F��Yw$�N��/ڂ�:��^�Y��[�:KM?\�\��^|R�h���#�]|ox|E�j�5	��/ת5!��luZs�S�gZ-�7�Ҍ�{�,$�ޱ+���HaDL��e����uc<�և�iO���\Ue4.0,���o���� �Ù5%M����ɧ�KvJ�jj��{��~���Ϝ� 0h�'�{A�m�tћP���V�����Ϻ Ə��=�ɚF_��CX����C�!����Y�v�^0<�x�iF(7�.S)�Eߔ��A7OZ��oUUtg)�5�i�����lQ����[�ZM3��鄺�z��۫��s<���Z��,�ADTE��UGǮ�����,����e8wB�=�m�Ñaퟍ���BH2�M�P`��<{2Z@��&���&�.�j�sW2����0��[(8��m��=+u�\f�I�q���:ΰ�/2S}��̭S����d^{���1����E�\�g�1#q��v����"�q����Gw�p��fK�ur|�0!�����+7�����Q�8��X$i-�W,�()��}\�}8\�D~�7����
%�����-dW�vW�D�?7
�%k0^P�k��swDh���:�B1����?��<oϮR���H�5@��:L4[��]���E�M�7�PPX;-�}��[0M��1)�u�`!�.��>��tx����ܤ��Rܐ���U�-(�C��ŗq;5m�dq��;álf�x]�o�?��|������U�����u�L��o�k��N�3�8TI������c��G��=?iر�)�F�dc�����\��O�E��c� /}���郓Cv�6���%T�=�=$�:4^����&�ip(㬸�=?J�c��"J���F�D�}�*�഼��V�`㯚��'w��='���k��x1�S�+t��%�Mcz1'>ʖ�I�6�Jɽm�8|���KT���q��\�f�(f[NhF"˹p}�.���}Pe\d�:D�"fw��kb1���^�n��3��gw�F���RDu��Sݖ^�/ϊ�&�LL�U��+��>Ci��1{1e�?F]o3b�w1X{�����n���FX�KO<�1K?�#�[� r���~&α1<+g�z\4tEn��t�E�I��w�H�7���x��<ګ�>98���N����\��)�Bw�@YyUp8X�Y����SK�3ǋ�"R�s�T�?���߼�D��u�=�)<�*�xv�[e�liD�/"n�� �0.I.[�<"6���0�t���sE��Jq⸘��[@`kP����>�ۣ^A����N��ɐ�1���9$�)c��Z��% �چh/����rh�hbLyH2h������W ��%�3�A��[����K����m�|m�Û�V Z�U��gC��cx��
��i���bjջ�J0n�{G3|����\`��z	k�jw�94Qٞ/S&�%����@0\��(pӏ%ָؔ;��P��	x�e�����+r@�/�+=a�)��u���.�E�#p��im��̂�/Ah��K\��{�w�N���<tt�fI妵�^�,��hPˍvD.���}
?��PͻA��1�%U���ii�ڱ~��e"]RxJ����W�.$-*�Ώd�����Vŝ)F��36`���2m*��2�����o����o�%i�s&/�\/G�hw딳���˱l��A�_�k������n��XE�@/�c��W�4�Y�Y�M��tX�����1p�gdO��Ct�r5� �p0��]:���?�E=d1&A:
�!�@åu^� �/���}T��Y�H�4��p =;c!6��+�x�j�i��><d�(<�}��f
$)�<5�!uS���{��L���wSv���&��b����¯26-�E-�BM��w�����{�Ň.	�V3����n�a��2�j�m͌T�A�İ �)�M�+oƭ��%7���� vX��48@��r�g��,���+��f��);3
C-6HZWWqrᑤ+]V��0�'�
I��R�Kl���)��8~��0�{�b��閰����QM+/w�H7S�a�)Dv��[Z��?�힖rՆ!�J��UՑ��a;���O�00]�xǘ
�����H���?2=�0\�F,��4����hVe�~wS	z>���,	.[ً4F姾�I���nmH3�k�.�*�˖MKF&����fY�hy����7� $Ϻ!�/Α��ӟ^����D�w��P*������ �\�}�4��[n~ ����O�[��9�A
�j[�ui�.M��M���3��]D"�)>-�q	"S����l�z������&k��Ι����17#M��IK�i�Qޛ�.P�`��j��G	�Om������{�4�9q*Q��W���oG��ӎ�g����N�7r���M3HhM���)�v���Rb��I�|�D��f�t�Ap�f�/�zD�Jxg�6�sC��X)5�4!����5�G��j��Z��m3�M{0�~?�l?S���>���[e��R�S�U���UPx�U8����L�I�+�	� �> �gRQfk8F�H�����x��Z�`m��Z{"�%@6�ȋo6����S[��f�򪁄 �����C� ����j��~���j�%A�I"��t��_-ͩ�4��� S� ��nѩ<\�'��kÏ}m���3�~�qjX��~4W�H�N�1ȗ%��8o�G}HI��  /)����:8S�XE����@���e/�*�a�X��V8-)�6T|����oSE%�?%�U�r<�E&�'$x"�� �����m��G҇������U󻁋#��1���$���	C�}��W���"������ ˵-!���������	����i�u�F| �6~��'�q>�[
}����
ձ@y؀���ϚR|�tw��I5�z��˨H��{P�U뱶��?e�3�ʂ�Bt@?��
�Ba��T���;8T��ӅG���RkߤJ�@z4δ4GSڿ�LÁ������bj3&���:���~7�BG�M�^!f3'���rr̍�'1���x�����O7'ۅAQ\��ރ�#j��΅�u�.�7�A/�f��O��eYۍMFnR�V���0�;$%��Zbӛ~���Q ���=����?���	89g�B0ϑ�;�c��
�x����fWZ�7�ϗ{��R0�b
����yt��Ř >�w���D��Z5dG+���f
�2ԧƒİ��{n���5�ڟ�h�J�O��eE����Q�R�P	X�x,<_}P�1�H �Y�;cβ��<��ݟWc3�"'�注�K�	��.b�K�������1�N��L��D��?,�zd����*,+l�p.�\�F�+�EeGK��x�5�96�d�.����f���(�����S;ʗ����n�ؾRʖ�~�H;0�=b����|Nm�&o��	�	a�
��g:(etd6�D�� [q��=�^�����%G��djKNV�����<\�$��,����B�B��l�`���o;2s=���n��|+D����'�Z��dɶR9��S湖-w;�5�%�K��V��[����*]��������89"Ӣ%]���#�[2��z��Lb���t���"w���