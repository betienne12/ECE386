XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����I�s5�i����`������:���3�����S��	~�"u�`j9W�<�ᘦnt�����U��?�*�wn�������J.��~�v���y�of����_Y�$�?'�~Y���O��rT# ;J�jy�iwu��q�)��qg��=k�3��&�L*���P�CZe3�6C�
��w8�d�]������i��$��a ��d�P���ò֝	�w�ʮ�89���;�N��Qdt��;5˺�i�/�T� ��}�W��w�6�Q%�JI�����hb;�qC=������+��}2����D��>��ɶ[��Ҟ��3�9;E�h�>�]�J�����L?<��.E\_�
֒,�Jk�r����Պ��j���ݙ��&�u�2�R�~�*�v���d����DXIݘQ8�"_�%-�ˣ�-�(q+.�C&���˱.�����q��{2f{ΈZ}�YH���!m�C�����P�nn�KV" Ӱ�m+Г�i�(c�����k���!�����!���D��j��)\�<�T��h	?�!��h.�k�t�p��U&�4o�D�P��J��F����:ǒ��:ҏ\����K�P'�˵�uH�8�����JK �sm���$@��c;��t>��7{sVں�kPz�@~��d&(j�e�{�{�t��,�c\�d��n�~�2�{�,���2�r���+e�����*[��ՆJ9�g�ᐨ�I'�����M(���e���)�љl���XlxVHYEB    7744    1780"�+�?aSje��=�\d����Rj�+�S��?�\+5A��,!�5�S�-v�"ɱY���6XCO�c�k�<�jU|��-=h��4�oc��S�q��&eX1*�4}�j\���E��8$��oo���p��=ތ����)���=��ȶ؃��֋;q�;�wRjZ�XR�Gw<64������݋8��p�A���C��z���vi��f�x��P"�Nm�NI��RR��x�z���Ol�4� rJ���51��k�飓���$��Ѐ����3���7j=�a�ר�[���bD��lI�f�ȃ/����`afi�s��-3�q\�$��xO ,���F�&^3�n�/O,m�<e�+Rc':�n�Չp�ZFi㺨�$��$�1i�}���ŴM�4��7Lg�����?T�Lם�pk��0H>��XY�sDE,�@��GK��q;LW�¾��9�&��x{,�/�0j��U�<C���s��ϬY���K�T_S%)��]��7��x`�!n�̡�,��J�R���va��yI�4#"W=���V���OM��p&b})����p�S�	�1z��/	���Qx�7��~�$@�*2�{+"�CF-Q*��*�ȯu�]���n3��ٴ�����;�^�r3P�FmO�G;�6fs�d�71_����W�*9���i��ui9�/� 'y�$�"����:g)��58�݅M\+�A1����Ь8T;Vgd`��fo� .�� ��&�:�5[]�r뾖^�M7�m��GC�p��Wk��~�����}�-.؟��_@7���?��RMr�:�a{
<(�^x.hm�K�����n��2��D�YJ�d|�gv�����#�Çk�V���u5m���e�b1��s��	T0{%�c�8�k��Ć^fI�]��Gm�P@�N!�=�/F�}�������Yy�x�1�'#����X�<�DE���%�9�H�
+-�(�,~2�@�v�7D�i�m�A�D���y�d	��Lې��hl��XPJo§�"�o"�Y����L�M����V��Z�GHj��Կy�D�gF�����	LG�W�_�г�T9�i�<)tݮڇ[�����L��\�7�[	��������`�i�'6��ޣ��Q�r?h�Ǧ.����J^��������=��͝O,�b��@V�߇c{���k�g34�s��j�Sf�Y���T8�|\ �S���͒k�y.�_��!�s2��\�`�������4���;i{
9,Wq�o=T�в���D���^i 7�(P��-����"D�C�F;4��bҌ�XvG1�Qi�`�0.��E��C���a�n�"���i����n&����{�7��d���� hP�Auy̬:?�����z�Sb"�:H���/� ;zڼ�L;��X`Q2j�~��>�E��bڠ���/�����'�!�};�Y(:,&T�s=�	V�6�/W@����!JB�؎j)������mn/�!XEec�Ga �'�^.��E	�/�����nٽi�λ��B$�%r�I�J���XXM�f���:�g����R�����ׁ(���3xLXI������=DJ��S�ɜI��	���7���'S��o$
�r��h��.; &�F���=[qta�*8@�<��a�9��:�V�/ �Mu6]�h�
a1䦺n��>sA Sl��yww�Z�3?rEo��i�W��6�?	�~1��s^�> �����X���M�/3f���!���t�"h#��Ǖ=���ll��K5�2O�-Mp�>>{�f���<�[��5B�N��  �!7">o	\S9�ru��y5�~�ބ �r��0��ܫ+�D�ͺ�L�݅%�42��v��	x������܅�g�o]��Wy/�Y�=�'�4�+�Z��/.c� ����D��>)�<ʴ��D�2w���{�*�G�L�ڦ����28���1m�^ñ�#v/��n�Q��rV����P6Y�&ˊ��#煲_',�����-)��5uTY�1F��r��2Z���xc]��aM	�aΩ���Z��#R!!�����y)q���~O�Ar9���A,:t*���LӤ��b����OZW�L)S4���3P=P	�T3O)ɭB� q�R�/���d�.��"!QZ�-���vf��׫�yт� U�d.��C⏓���
]�=Irn�p����D���,�V�?�<�S��m9Z���b���oZ ����X��J�t� ��o�z`��U������ߤ`@	EXȓj? �X�ȩAM@P�g_��o-p,�ʸ�m.{���<���,-��fnt9��h�@�\m��.��
�Y)2`����OB.�ts����Oum��JkC`5d�&��"�*��k� ����{�Bn�0�ۅ7(/�%	<@�������Ͷ.p�Y?�%-�Wv��Xm�o@4���."��灧r�K�-�ʵٺk:�a�
��\e���~��$B3`��_�����#���f�+���[bnSq;�Y����ó�BH�'U��sٶ���n\����p�_���z��u_��ݔ���,�B�#Xʥ����Ί;��٣v�HBk���S��A�O����tg�x��KK�SҖ��Sf}I���o�)��@B����]�=tuQ<�M@D7@t����?�{X��V_��C4�-*! 
��h��?����l�e��D��A#�wY����i���e>1�2@��8A�
��#��YG�2�,�>/�^��lC��"k�����|�p��#W����8&1����ae"���q[� Ǚ'7��[�� z��|MH�3�_������Jٖ�:�##D<���Mt!��@M�*��s��
CS��;un�g��V�q��& ��R����o�մ�,���sl���L�j�ˋU�6'��W1�a��]��,Z�;��Yj�I'(��[�^Ld�eJ`����[��X�n鮗�Đ�˴��Px��^��t,�A= uF�ߏZ�5�|��|Z�d�7�����N����G���Und!��(�J_|Z潨1����g$��h����AD��>�٘k�n��I�Ń��d`9�aC���R������9���T�λ�"d̒�0���EZ���\� ��4��_��f� �pY_X���o���!+Jk  �:�pL������G��bŔW��+A>f>�x�mഃB���R���P�$h�=���^��݂ە�j��|x�"/$�ꭻ�#�W�fB�.ʍ���!=�'"m�8�U�#7�#M?�Z9ϸ0���i���:ޘw�L���H�m�qc�9~%Y�#�����,��ߒt�O}��\㌹}������+� 7g�����<FM0Z*�����ȫw��If�m��%��8�|s��/��ߟ;c^�:����(��������עiï��q0Z?����Ie�!�q��o�����&��[�d@1�F�:���^�I�����?k��i]k� @&�/*�k��Q���	)���̽�Tvr��ψ�szg���]�ԛ)!}6����[ik�R
�A���p�ʗH���1�2=k����3�Ȃ����������*@��k�?{TT�8���@��?El��1A5%�_ ��S�S�.U?X��hy�z�ݦ�>TCj�eBڱnuR�߇�Wۙ4&������פp����S�_�?�?��n&�VX�����N��h��	H! �Ƭo��tp0&:���u� T���3����ul��������Dڤ�>Q>�'����T�8>���h������(��AJ}h�B���s�#G]����'E�`����="( ���a����_q�zW9[�<�;�-�/����&�᧽����ZŘ�bMI�Z��*f��!|3 m/��f&E�}j�H�3ZIU�4"W�}�qG ͥ�$7��>7�<��G����-��FK������V�"��0��Ma����7�VJj�4�?).�iX=���MW�ߥ?W_�^�����ω�V���9�|y2��Z�?L�!]��7aK��[���*@����]�Z!BG����󵡕�5LJ�w.����2
��G������.5v%����N8�x�?�F�F,���v�,l.̠Ng�K�rS�2�٣��^�sAf�e{�W�:�ԍĖ�OӖa������5�I�5W�#��A�1�Kq�5�%�]����:�K(��mV���<�$3m�a�& U���L1�!�ƌ�-~�e����3�R-�a�����^�9��B�z�f��}V$7�� m.�	<E�
�j9o� �z�ښ�C[�C/�o� ���2	����?Uv�L��������*��_�MV{+=KZ,٦S���}�R�x��d����"�qEUn	C3Cx�Vh޾=�hP?V�+c�A7�@���+!R�ڪPd�C'h��>�k����Ϋj�����X�O�u����<� ��P����qb.�紺�}_ | �c���@�_+�OĹ�Q�C'0n%�
�KO[�@ةQ`]$�1 ��"���=DR�X&�	c�RSS&?dr��5�@;���܎��<B6z�ݰ2X������=�p����Q��Q.���J)���Y�UbTF�[������^D�f�"yjb>����moo�8�M����.�ėF����,)䣍t���㟖��r��,�E�`$�A�w�W�_Vc�~��:<M�W�Nڶ�9#��ü�KnB��6��h���T�/Yx&SMPA���e�
���o��_���,�6���?�$�vl3cN%�:���X�^raIE�<�e� 2�Th�(1�����tX�c5p��(�]�Z��������#Y��Xhށ�'�����%���wjQbې�c��/�ᇳ�ƃ0玚,�(�G���-LN!I����o!Ft�.��PF9�D%b4q�\�ŭd�yD���H��)._�;����>�:7ۮ^���)�g�Qz�&M}J�[�;Q�������=�d�����`��?O�]��2��(�?b��ֲV�8*̑.�A��mQK�Z�j��x:��8��"�-��S8�A��������ً���m�r|�A�@sC��"i�YRrR���Af��s%H��hV@���L����@���/!��
�+����F=?\�>�P�ზ���`���H��T.��q#�^��.�@�X׎)�^���{��l.���i�(�m@5��h�BI�k��5�����C%��S����;��>R?h�-���[��.9��keRO�Ӏy�$�q	kp�ň+�A��������C�>��5�j#�����E�t�=���h�����|_��4�~ �f%�ԗ���AS�~���%+E�h��䎼E�e���y��	݊&�	��Z1C�#2q��|%!�֔��Ok��'I�2|�#���r�/������!��o�w���)�:�/�"���J����F����6kz�Hא��6pU�`�n˟Us�~�|ϖ,��f�h��y���zˬ�J�xE>>�.DM�R̝�O��*R|	���mUG4����#�s��_2�y�� ��%�Jv���z����K<ϋ�����D����!�_���9[�_����}Q���b�.|��',Kw��� xX�֟{��>o�B3��Y��!�ɫ�*lĥ�S���C(�*BO�h� �aR�iq�8�N���$��N�]�����΀��~�[���N,��7�:s��-�-��t!\���KK����Ɇe$�=g,T�غF��7�p���S�Y����N����R�jO'�k�^�K"�;�Ej����[�_����r�j����z%+�o��6$��s�����1Y}
G�+s�����N.6��V�)���*;�4u�V����B�y�g�O�c��5V��*Da'�pq�,4�leZw%A�i��h���v�l�&���S�L�