XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�'�WrL^�࠯��XseR�,%�l&����z�
rٝ�����X���ѧ���5:��lQ��e�����?���n)Te
����d���(U�b�@�x�7O����J/X�{e`�nݨ�R�Դ1�k9�BR�}��+��	��;	
�?@�1���L�b��K��b�A¯��5��s�%�u���zs2��_[�dȸ�|;+�~�x_��b.��ԟ�����tkj�3�����cp*[)�b]j��μJ�L�[:U�E� L�)1g�Hu��]�sc�e<u�%U�m�N��⦦��Sf^�����L���:obZ��љԜ�����bK�A_���S�gw6�vt�0Zj-��0�����`A�pڏN!���1�����SDT�U�d��A�9��T+o�
�M��;��"�	�xC��Z�$7��?�����ׇ"�M��m�Վ��{���,kh:��r��&��P���i�C��<z�DR/LVH|�.�����PހV�clT�kc(*Ju.[�/��b���2~��n�얐(n�)R����)������.�#t��
J	̂��� c��.��5�+�*�(��#��"�'��p~���]�%�
������B}�dh�I1!�S�S�'�w`��l�1ɍ�dW�{���O%�UIu�9����x�!��/�3!C)2X�vbȽ{�nD��/����U�.�D����P�T0�םlP�� ?|w��#\�ZaG���v���na�P�U��z�K���vb��;#b�W%�XlxVHYEB    c763    2600Ŵ�_�V%���{)`SP���<L~R�)%��|����iz��~��.=D$ݤ�C� ��&�C绚4�I+��H����^�v4Hw&�"��P��>�+��в��wX
g�n�O0��ujߋ<��|�%��Žǧ��˒�u�hk�K�ء���rۭ+y��@!�b[H�������(�`�f�~%)����fۑ3�n�9#}�_�e3U+���A&�"QD�I�(��%��Z������]�Ϭ�G	�'��ii�ح�h�f����{��Un�P��7q�D�Uk!2'�%!���������)-#�:AI�|�;7`>�Pʓf�4RrGhk����Dk?�.��|@�01����[�^�d��2a��B��8��<�0��XD�� �҆��Q�Zrrݦy�DI_	��#vO��\���ͩ�
����W�F9b3�6������oe��xJvmwr�x#Qߪ�Y���/�U@���|c�������?�q���i��M�ctAT������+QZ��0���Mƃs�팴>0;�h!$��img����S�乳?�5l�!��A������bb�_�QЦQ�=�� y)�]Z&a�C΂������B^F?�ю�&5B��!����I)F���W���fv<�S�iKE�S�N}����r��)B���ۥ�Ǒ�7�F��h�l$�r�r���5�<Ƞ]���'��(83���;��)���D3��l��.Q�K@���,(�I�R�ߢΘ�jQlW%r�+��v��(|<��T���&4S��/�?��>e�p�i�:�� ��2"�hw�4'�D�A�	ن0B�;?ܕ�)�����z��A���~J��1EQ��Cu%�����ܟzܓ�u����0���x���B3ޚ'�� ��k�����wbw�\"E���p��)�p���������!I���� ��ܛQqH���"��}�/��[���r0�K�_&��aҚ�c^�����O�j�i�/#�YP�=)ҭ��P��J�p5�/.��<.���.
�Y�b�~�a�!��WI-���	K� �2*�sᏑ8|�^$�V�y�ȼ;szI�o�a�Eެ�Ό��}?��*��'6�>��a�DG._M���;�o��%��%�Wp)8��4���݉�o����W��QB,^����c���a���gs�7�F�@��qug����}����0�e�vr�� �"���l�ZY3f�s�)Bh&�`�"G'�) �G�)o_��,�%h-�v��<�O�R�FM�]6۫�Ћ�p!	�9SC?B��we�!��ǖ*У�\o��"bU�9�2x7��Ѷl�F`�#_h�����W=�֨24�`�P��A��#�I�����b%��=��A��T��w��8���!��ou���P>O!�w�z��=;��R�+@�5{Ѣ������JIj�u��:Y��� ��?�`l�Fv��*�����m�J�WR5I����?�h���~�L�����~�=��qqq�z�p���k���&���_�q��Bnyj�a;b��kH�,ծ��CL�]秫��ްr��k̬	c�E��v�͹G�OC{���'���`��l.��7��M�K����,���p}'ۣ�K�GTZ�zj��	�L��H����9��*F�í�d���ϹQh���8Nfq�k�0f�?ހ�"0բ�!�f3���(A}:�7���U�^����班"�y����$o�দ������:4�k�C��Zx�$O�d6�� $�v�h$`��e:D���c�3�&��F�5����rl��ſ����^��ią��3�X�>H�-qI�����$�jAj�9	N���y����1ș�$��X�<0�-��t4�u"�BM��v�ˢ�`5u��X���[����������� #L�r+=�źK'�S"���B�����#��Y�q'"�4�9([ً�äO�i:Zŷu��A���ʔ	�i�~���I2��>�������g���r!�z�:X�0}?8I�ns�,B�!v@2�~��qɗ�+j��K�9)`�D"g��O_+܉N`]X���@�������mm�wQ����%յںaL���hG���n���{3�[٭�ߞ�q��8�s��/��=&��D_zXUwB+u�)��/����w�	m���n���#穔��Ѵ�����
H��-\�^}�߭y{2����ņ5{�;a��4.�Gc�ᕒm�J�}8�O�4��/T��K�ѐ���_T��D_�W*��i%��Эn�����L���t��XP8]5�a�V-h
� |���u8��ΒL��kr��V��h����zw�Yɇ�Px'
���u�2�e���0�P����vd�փc�0�����L]��V?�@gUW�3]Ӂ�B�t��w��pO���}N��'3F��_��[pN�j��f��W�)�.���y0a�Ua�F	�G�O��@t%��T���#%�[�?F-��}�v{U�=�PE�����h�������g�>�$.ޚ��o��u�v�,��~*(E��;t�O;��E�Ndj�N���h6�諂�-��B����v(��(FW�W˂���[
J�������,:�Y�qn_{ ��SU'��#���WxWǅ��}�?�M�蝝����������E�&6Ft����)�HD�]��R���d�{�a0Ņ�i]�P6BI0�)�Q�g��܃)�N�P�2�&WeN�3���|Q�A:9�.�I �TNP��j
1
"�����]х,�'s�����I���Ѯ��!@`TS���o�����5�χ>��ʹ�j($��M�#ŗ�2�:�b��e|ʌ�B ��KWve�~��qZ)Vq\�׳�\m��}��8�\c/7�� Sk�j��s�/]I��6���=�2t�Pߨ�C�}�X"�ۦxZ��k�rfVH�����Tb�J6Bv��m��T�#AdG�����-c~�1�+^���Y��u`ց-��-Gi���k+dv��E�e�k� � �/v�S�EiI��m6M,�����4�ђJ��J.ގ3m�yz�㐍\�ρ�H���c��fݥ��w�tC��6�|I`@�T����u����F��B5�\�K'6G�����U��+�=���@��A�}��M��p�;����&��G��]�N{V80u�;�2{��aٰ!���!A�HS>Z���=(��uX�gG�)���Q�V; ��|�
�Gk�W+�w� n0Q���?�x��Z���=f�dp 9*���T&0<�Ț^Zt���|�� R��j�,��"�Vh|���ܨ�����@Z����ߩo�<��s���3�u��?X铛������ 6r*,E(�]4�S[[�Ec��(P�j	,�G�;�G�ST����	-|א6?j!M̏^�u�������q%zDBN�S�&��SC�~���?�ԭ�`lE���[y�����%x�hqə�� w?~���*bf�K:�嶤��+K}=w�o��f3��eU�m�o:%#�4�+
�^Js�]p��٦�nc�9����ʄ���m��_s���&x�7�wc�� ��&�t�)zHH1b��w�n`M�z�!�0J�\���Y�nT��E�밁�&������v�ck�h�o�ڒ8rB>�>�T���m�~_�IX����eӓ�u�+EW�8t�[�#S܄���S�l'e�2[!���Uؽ�����h��]��K���ٮt
{�@��^�H5�yLȩ�)�������^�#j�ĮE���D/f!�m������,c��r���ӿ�۸`w6骷Nm�}��x.���n6����M��T�T�hc�9��<��]C��B�p�FW(B�Sa��Âu�3�u�,��mĸv��Mu���q�e'�����@�.?�Z1{�]o��}J㒲��g�孂�/(���g׽f��E��6�Z����tm��Z��(X���T9��R���go����e�>���?3s�F�Vx}Z�m�Y-j�8|���]]2;d���ENv�ϖ*jJ	M�i���z]w"�XP!���'���l��}RiO�%$}�5]���$���W�Q���z���stdC���ĉr�n�x�G�Q�]��#U<�Ļ.�g�I :b6ޤ�9�>��گ4��sʯLL�u1)X�7[J�j�hrJ�x#E���r/(�)|D�_\]��h�7�����:�]����!V1����Ǩ]Z���~����EC!�w[��G�3}�]�����E,�v7$O��&��6���h�#����U�R.�zl�=�P��j����ܡ���OA��#rj���E����#7R�������zB��Xk����};0�(Y���R0�gi<ڨr+��)�,U����e&$Ⱦ�i�\�4Z��U�%�}��%�us����P	�X��g���Co��FhB7�R�OJ+t�)�蝊n���>�b��\5���b�8f�Rj����CB�z����`�t���%�^EL��aWQ��]�y�f���+R%����\~���z��"�����q��gh���"#�@�q�?�2� �d9#�71t����K������#*�rK����A($� $��m��X26�!�|-�5+��f��씋(��2uCL��܉��>Űw 2����c��@CŘ"�l���G�7��j-�T"�-֒��hv�*��od�h%�C��R�+$F��w��;޽�Np�'r��Gbi2>	�XB���O\��@J���lR.Qc�y4��3�4�����1�>�r�R�w"e`-���9_��fdA�aQ2���F ��ԖRn��
�s�k%��5���&���;����m����I"~�3�S8�
���-���8�4�~����NԂ��	mx�1�"��b�I ��|��`��&�^4g+������E]hil����:��p8<z��h��YP�������J�)#�` q5���|c#j���?q~h�u}�Iܱ��P)�������DJs�_c	R[X���ЩJt5<��\�c���6��DdbO�)��ӛS��ʽ�N̳?y��ڪMR�">#D �>Ǿ�8��Wʨ�{�n_�8�ai��R.0s�J1c	�@.�qu_��EX�G����)�(C������\~g�&�ۭ�����s�P���D���p�1�4���%&B�%��Z(�5ڂ����X� ���ȳ|�vt���CX�u��Yyb�R���'�e��)@�~8V�7�+
�-���u[7��4 ��\�.o�AǦ76���$q��TE��0�|��i-l-qy�Pk �vCm������� =��:�Ӧ�Vx3����M_'ĵK�pr��3 W��0��_b#�W��s+k�2�=8_����:�QK$1t	1M ��&�nC#�(�u�V����p	pm��1W�p��⩤�[e#��z��$����A�
�������q�(��P��9����B���09���n%fN���D��I�^W�y��&�����.0����ʻZU ^EW��,�s B��g�'�����m��r�p��u�hi�r3\(��鐲�G�� y�z�b�6󾻄�����{J�lKCa�1�����P3s��n�ut!|��l�֊�vw� ���fDY�9�����+8�3C��*��+���9@�֍u�^}�
�њ[�K'��׀G`P�ۼ��T\�6[Kz��J]&�e7�;B��B��-k Ƅ��p�.�8cQ� �����Yz [�Rr
)K���?�X�ߥ���̆�W��σ���������HC����e�i��8
�~l�q����4��#x����-����Q%.!�i�Y�qt3@�#È2Ġ|��$�ֈ�;�����2��do�U���Ye`�Aks�r)�L�]�p���Y�v+R1���>�g�;��J�U١
���O)���P���l�EV�%I��j�x�54��\5һn����[:�qs*�.�|�˥���;Rwq�<��g�b�R@��a�X��Q�� ;wŪMT��6�%+��#�1$>q����7��D��lG+�g�8��О��J���{��=C)n��P�7F3l����)�qn�Ox���p	0͉��ۢP�LC_.��d�gG�-nC�8۠�A��\��&_�	�R{�����U�唟V� �m~�+�~�ʇ���	G��?���xNz��#m�,���$�]P���J�J���V�q�	��`�e�W�5���}͚�W�t���Qi��+j��ᗐ1�-]�Ϡ�����������'��>Z����Y^���T��;$���I�Ҩ�:�{�'y����%c��T��� y�h�
�G�\�����L�Ж�b(���.�����NX���½�'�$���nO��w	���$�NX�1�n���O@(w�
�N��\|����+���3���� ���3��F.J��8.�F���ǘ��)E�t�Ɨ��ޱxo:Զ�z� �ö���~#�.��gކ��>��Ɛ�̋��C�����<���clݰ��:�1V�HI���Az�)��w����k98Q�7C8@$*�`��C��s��;E5�ˇJ��UWL��9^���
��F����G��\����4Ѥj
�(b�&K���0��ثvUH�$�~ה+w+��慁��_e0ϖ?�b�Sr^�3f%�����2{p�U^K�C��#%v%�� Ɠ�����rB�>��y����nXi����CbƫfS�������r�0�.*�Y�| 0��	�Q(�;��0�w{��.���YGj�iy���$Ta��|���~���J.�	U����b��D���<����w��Z�V��a}�f
��}��NpTU{�^Ifz6��2�:&G!�R��VS�RF?�#�G(�>T:��H�O�k�����Z�_����^aJn�/A)�p�l����M/Wf�L���Έ 0&j�e�}Yة@T 3�V��=gT�,�� �3�[�2��!��t�ʼ��~^�Ѥ���2�+#��>�`4Z5�\v�F�6�Oޛ�k�m@F��Mfۋ彯u�Z�Qsv�57/��b���i^3�j{�F���%��LTح¥�~��jȭv7�%VGڋ�6e��/8�L���M��=Z�5wO�L�JGg��>
��<-�����V%�X���\)Z�>�=§�P	C(�Ɂ�L./������$Y���
���^���6/�Uߵ�~J?����y�,�d���:(�ɾB�˦^�hZkf��5���
�$,g"kLY�/Eq;�k`���C_b���g���T2�������"ӯ!Q5+3��yj��eD�jb��N�N�bM(���x[��l��D����[��u�/~HL�C~�@�QڐTK�aY�f�A�� ����d���p+/�p����������-@ y���ug,N$I͂�|`3�{ 8�����$kF�Q*3�����U�d��]wz��.流T�M�{o�(��*�n$M�ժ#_�-������ó���&м@&��?��|�G�g�R������&�������Ԏ��%��E_�qj���b���W3�eVO9�ꜵD�7Eҷ���~螜 2t��5�Z���M:K�7�Z*�#���רs���~��%{��'��n,���fl�80=dc���WqB�t�#2��Iƺ�\���j��'�X�vO&T�dʥ�f�gϷ^�a�7s~�����'�n��P�lYN�u��7��g������kz5��H���O� C� ��4�����]LH�*��.yWu��Q�
�i�`�A�LL���]d�v�l �� J��^��N��LT��rԹ�hj��\E�h(]���t�6�I�� I�#�u��]�3 ��Q����R���%s�v�J|~Ex��$�'�]�NM��������ZR�g��p��zt�?��M��C�"� ���XS6���	$�Q��g{��gX$��>�͇F���2����8���Ues;��\�Ai�|�Tê���>'4l�)���~�Y���EK�;���o�GE4_��P�g,4;W`ˤ`,�Ɲ�~�RpW;�T�3LS��q��
x|��Q��_}i�pS��S#n,�Zq��B�p��
������DZ�K�V?y��>�U���}� ݏM�x2lO�Qs%.!�I\I���!j���~�9^ʋ�kwƮ�~�-J��%"F��pq��6=�U�h`+��A�A� ���9�q���f8�{�������+)�\L���?� �
���beU���4j��},O��������y����BJYV]m��
u�&��ˎc����0���qQ��c�W�0C���ms��ۜ%�2�s'`p-�\����#��]`-�O���3�*'w�g*GV�:����ę ����:��X�Y{��� 4�$9@�Aq8��EDǝb��p�PД� ���8/L�B��p4�=E��P��թieȍ׷�~�n�10��OF�a� >����w�g7�D:uxG�7�za:���;��6Lr��]��>���IX�j���$��{�ژ�H�e�֭�
Wo�B.P�!����tm�\���/�Fk9�`�1��vdTHby���J���DsO׵���iƮ� `_DZ�O�v�S�Q�\��\��Ek`I�ⲅ#Φ�1W|x1��9��Ѡ�Y�}D?j����98�R���^�3g���r�C Q~�T��G�x����kUsRO���a�@.QNZ0޶�������s��1�T�q/��|�i\�3��ڱaEF� �s�-��bk���g��|��(�T���/��ǉ[��Z�S���`���R&�A�6a�j����JHe�Eq��' >�x ��Nt��#9i(Y9S((43���9� ��V3�e�0c1]���F��u����2�'G�І��@����]�:V|樅�f=���|e	����d�n��l'M���<�u�q�%͢�΄i���ڽ��ǒb2�C��#]E�=Ӹ�'� �O=K���a^��n/���1�)jZ��మ!�Y854���nIyoz^v�	�{�!鱿�/���1Ņ.�n�c�4R�@P��p��q��������:w*96���W+8�D����-��#9j�FʘbN�r�+�[���	7�?�#�������|��f?}��y��V����2m���y4�>[r ��#͛Nh�����aj*���N�eZK$�>L�kO�IJ�p0�����GK-�s�����T���Q����/ �-����
�Z!f�Mo��u_%<�zE�TR7���縕�G����� ʰ��"�����Ϡ�,)���#
���]-B"\�|���ƻ�:1�䲾o�t$yߡ��av9�~M2��"��w�%h}�����$����k��d��Ť��t�H��q�FK�I��� ������Ϻ�n1c�b���)��"��1��+�P*a�E��1�y��C%�E2��\7$SI!��BSݦ��<