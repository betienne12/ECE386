XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-���yN �=��� ���;]u4���ޫ�`�����
h�Q�Qq�}&Z�qeɴ
�҆�x�i� �2���<�10J���4��)��5M�����<1������|�Rl�X�(D(���9�����)��E�xH���7k��tȂ/N܍:���?�Z��#݇]�|w�EX��1$�<V��Z[:Z���np�ӰAi�N�]a����T=���̾��1�9s�;�>��]�)\����R�p���u�̹ 2���PAs]�D@���T�s	l��jp�e�P��|G}���AԜ},k�A�	FR��Z�dQn@;_�b��y<~�T��Y�V!<}S�8����L�C���P�W��&lA
=mn���>��	�{&�>��p����������������1{�F p�xZ��<	��h S#���\���P�TR�V�:D4�������;z�:f�&�ε�Z��ox���L����a���=�cx�G���z���ªG�m
��^��q.��-P�����ޙ����V�?[[(�o�N���%��$qKf�ׅ$z�����"��6�d�"B�%a�i�,r"�jP����cʥ>�Х>'�Q=|��a�j0�(
V�7Y���ŉ"
�����l�n�>���vq��ݑ҉G�iX���`�gs��[�D~8� �X������Ï��,�R�G)Z0Q��uݻ��SK֎��ݱ�$zi��! �?'Ev�#�xǴ��]s���$��2���XlxVHYEB    fa00    2030�@Gߜ���)S+�DH16��O��;���jDAx/�|��8\��W�f�>�D�M��$���v�7\�đ�� ���ڭiz��ࢵ�Su`�^V&)[�z��d���Ub5�R7my��5���˹�K~�`�y�ob�)1�b�߽���4|jkm\�|t��1�z��7)�jı3�`��d�& �[�~���ԙOѰ�Zm���T*��B�K�8rq0Xe�p�/��������}2wqNl�;��?�u�ą"(�Dh3M��\��~��W��J.� ��a�I�W��5�{T�1��D�B8�%q��@��2�P��>n=��lT��a~h����p���	�5���dj|c����ĭ��0%��,����ۄQ��5���U��x��Lf
�9���f`:�+գ�Y����A�١/��Ě�X9����츎�̢M��O2�1�o��r��p���v�����)����;?�fJ��B�Eo#\}�	��9W#��=�A�%[?%���N���Rk�7�_�s`�E�%\�ka+�w�v{�A+;~��9䁧P3�qgS~W ��~L 	�$w�Qڎo�@�}]�X���ﻹPf�5�1"�Az�������H�3�<4��sE�m ĝ�������h��y�Ep� �kϬ����G��fK ��Z�Z`!j�c�v�A��"w
�E�����L�� �T%*]���{��R#��:,I�ݍ��*ӢluO���2@�L í�4@*�e d�]� ���H�ǥf��Y��&a��=Oׁ�����#��f�ȏ{1F�R�N��b���	�*s��Qv�o;������H�T�����;��˾~T�n��!Я5��nqܽ��z�O>.c_ H"0���ʊr�-D6��3��̀Uv�J��O��,i��9Y?3Ϋ���Oؽ�;���(��۩ƃ��[LI�  c��,߁'Pd��;2Q��Փ�$��Ɂ�!�(9��G#`s�����:5�r�Z��c��b�|U|��~]�Z��G��4I�U�"G����uD����1��1�QH�Tz��~)W�qe�Y���#�+�B ����￼ڡ����<��z���fB�6ㄷ��5�謜���k�@�������#!i	��[�nf�sZfG�WrȐ�9E����y���P:��4��j8������|�D�=����4�T{è1��֑{R�������z�-�����J��i���*9Y�hw�� n��Z�a��������4$`��,�Դ�\(R�n���%�UB��*b��Z�ri���~���-�WK�]�g#8ݫP?���Il��k�>>O�2��iɭ�f���J��7��)�41��YT��i��tˌ���� \Z����� ��e�8�Cd�/��wE�rrx�4c�������-Zo����@����C��R�;���%G�U>�])J@O
�\�
�C=O����qZ�2<�Ê�ޝ�w���f_ �倃�k�����Ub]o�mH��t�^�H2'�O��~H�n�����<6L/��`��z�kݕ3����sI	B���\U�+pW�O�=�fd
y�@J'LY!ּk�*�.��F�Խ$��Ɓ��p,Z�z��>��ם�#�ߔ��������6��z��R'���d�@v��t�i.E�W��D��i�a�}`�#ٖ��7)���]V��ఽD��{��Wm������p����%)���|�^.�X|�k*Ӂ�(_
�����6�cPO�Kmz�x05O60��7��я�	K�=��O�aF'n/��
�NqIL�-5����o�J6��br\K2o
k�$�=۸�;��m^(��q��h�ȯҶ��eERl)#j�nFF���l��D�>���#J?��=�F�:�#*����z�2��9N��*�8��T1�p����K�C.8q���	�N��O�{[I�/��6��"�$l�\��Z��佬`��D���c�jȚ�l>S���b}���b�((	}?��U�n�窉j\BJʮ*c��)�y��%!���`�SRj�]�Os����8��!o�	���}h7O�-�Ƒ	Ű	�Ո�"̵39��u����sԑ7AI�(~g��~r�� t���l@�Q��ظB��Bx����nnCx��vD�%џ���kQ}h��n���Gl����U6�6�x����4j`"m�`�5����$�
��M���f��Px:%r��>�"���L@o�p�o�x���p��.��v u���S�C�c��Pv���:�}D��C�.Ra�����_��6ֈ+��y9�C � D�����H`�U�i����B�yN?���i$5�F�T����j��4$�[z5p���.M�4�S���z$���O$�g1a���)o��^<��i��^b<��<KE<�ψLO�T����H�A��@��Uzla;�xɰ����1l��ۚ�fS3W�<�i���w
RZ��>�p���� GȧqC9P�j���UᯒB�;����[=��ɠ�Oa��d��u����4��֬^h��I�P�ዃ�<U"�Ag��X����q�x�j��� ���F��wך�e(�.�3 ���E2�=��U���X�#-ۦHb����~�_w�=
��2�����!3��O�&f�!W���ctZ�( �!�5�e?�-_1N�$��n"L��{����������7!�EU��@��(����Q\���#:����+h#Lq)�� %E�[k�"�5X��e��e�8ɾ^�4F,=H�y�ΪqH��`˿P�f��b�p�m"�ek)�`6����.$�������_��n���S�`��U�%̰�؉Z�2>��F���6�&�K�S����[K\�bĆ�Vvos��R���h@mŰ�6�
m_��8�9�����j��u#m,���&f�4��������� ��RV��h���Gqc�ٚ��;פe���K4�>Á�M�]K ��Q����%���UI�W%��I�����$;�4��涼�pM��������
��&!-�0��yR��Z�2�	��e�[� ��!? �A�ȉ%�p3�� V0�=:C�RA��N�}�gu�t
i=7�xa��9E{��4�I��|��U]��?�����P��q�9f�əʑ�ٰv�[M����]�he�U$�%��І+��e�#{��7�ZH��~�>m�Ȼ'���� z�	X|\�rxg�b0�Bv-�Wl����D�&��gd 8�m2C���ٴ^�����잮s.�����{w�h(��� D�;OG���}��j\l�@���R�)���UF���[�lE�z2E�J�Y���ɤ{�$�
��Y���H��
rb8z$���6R|BQC�o��4
�˾'_�����hljأ�����N`�����~Lj��o	�5�.R�2p`��d�z�m�#�q"6 ��i6��<k�&�:Dq�]�x�a]?�n�7Ch�ϳл�N�o� l��_�lÃT��n� 	�M��Nʡ���>;��K���ҕ�|<�5�0S���}��.����&
��}��*�u��%	4D���T"F��O�档8 ����G ,Bؠ���{�:��+��X�#6�2�C�Xm�]�
i�b���t���~�[����s��?�c�Kb�[��������0{v�lo�s>������ߨsGx��\��3�[�,Zw�`�@/��l�&��Jg�xD�B�l��x�5���9B��;i��J���j�L�Y`���r8CR��v��N^T��� ��>i�Y�sNS�h�]��ՇcZ��?
���M,�Z�S>�-�V�(�W�PI?�(��2?�_�IW�Y�W���Mc�ۆK���e������I`p���e��vT�韬\�9���[��?�NZˉ��ҕ�&��Ԃ'^�l0�F֗���۪eg�HS���,!���a���]-5E��B�N��� cG��� d��#?��0����|:w���t�,��[�[�����2쁔�$\Yx��)����N���l�l�_�Q9��M'{��D)�f��C7��h�ќ�\c1
:����E�����Hk>��Ly�h�"y�u)��sB'?ɚm`�w����P
�m-��\:���B��LT�'���T�A!�8�� �4n9�k�e�6�)O����9V$7$I#�S�7*{�5K�"Jɟ��H�Z�^Cp!��q[O�V����{hE���2Ӂ� ;R4/�ਤM��RŹ][)'�n�f���1���kw� �,���D{\�YVh�������	=?^a�Dg��V`�XC�u�LWo��E6�>�X��+�ނA��7q�kOB3�Vկ��9���m،�F�za��
�i����z�6�.���(-���ȝ�_���#�_a
��w���T�����������-������0t�e0Z���sڊ�e��aS�1�%�y+������@�EI�@��q�	�˪��Y���	�M(4i�ۖw��I��^��_E]��7�K��հKb���~�#��{Mʙ�!��]&ڶ }�������6MJ�ۓ�z��/D_S?��f����lf[��C�r�U��i�?֬?�5ŋ����J���5�G�>��(]V�F]�����H�)���"~W����b�L���nB0�ր��g�>+7c��F���^���!�Zx]3�醁N���K���v�y��.X-��O-R�:�v��,���sЖW��X����"v�6~$&2%�T$!�s��5,�FSl���o�Ƿw`�u�[��bX|4=��s�qR��#�X��sW�<V@�%"f'&�(�|�'w��,�d	�&=U0R�"nN��	�)��~�1���؛�^���I?�gn$P�=G���_ђ#v�^�/��.��.l^7MR�le�0�Ι��"]�D/ɡ��L���ZgzB��)3]HkՌc���/�r���TW��WV��+��ٳ������P��&�������4ջN[����+8�����P	i�x�ڏ4k�j8��v�0�ϕ����{�Ǎ��%}��V���+K	�Km�4�Ol��%
B���YLA�̵�5$�ᖂ�W�_lT_����D&�+�MI�U��y��
D	S��%k+A��[|%��&����ѣW�������1-*ı�]��Q��(�Bf�Z4y}�T4���ܰ_�*6 '��yZAu�*Jј����h��w�H=�@����\�q68gq���2�]�N ��\�}źEn�q�ˁX�����B#��Xv~���:��H����^�e!�_�1�M�g���K)�,�T���y&h�s|���l�@�]F���23�.L�����ۤ+(��W��X���W��詝���Z�8A��X"�<� �t�y�b�*��<(�c���%;]H��Z�	��X_.-�
�o?~�En䶿��K�ȩ��ר��"{�2�>��]�\�rB�������5-��Y0��I���z�\ň��w�V�@�T��~��ݧ�|��c2�[��NcHB�� ��r자��F��~�mSR.[x(�g4�G+�-�E@T7� L��eˉ����[��.����\��jw,���uG�b�Z��o����%�jE���r9a�J�(��m��t{�%v���s�Ie,0A�^���g�/���D�7���0lC"���iHe���h��v`��G#?il�?������о93H���;�M1C�;&v��y~t��Qo���Ú?�Y�t]}�e��m�zXNItz���ڌ�9I!?r�!����m�V�,��(�3����=�q�!����
������+;��8��Ǎ�d�B�բ����?�c?��̴2.A�x�/�^���2��^�|%����b�C�:��<~D�Y��.���kF�>���i+�l�>�h�.�_�����;�)앍y�1pD�*���Yᾞaa��s��oyO)cF�l��JP��/�Yp"h��������W�9��G8d��B��PtG�'���h�#,C}�z��L�y+`6ds��up�Rl�����KYӥw�y�G�p�mC\,���buuǻӔP0j��������=�G؟+�L�U4���� (�DЧ�3e�Q��u[�C�0~ï�g���7&�y=��F��6r�*3~�ًE����޸Q�jƐ1�6߄Q��#��N���`�4��P'-�!�j�?��SI1e?��U�m�l��L�������(�]�?B�Pdq��;[M��y���}��N�Յ�6,���cĽ,�3�Y�OF0y@�dG�F�͌�g��&�& ���T�� ��A�46"�f�G�V�6TS"J�K8��0�i\���aά��W?���9(���&x�x�J��+�?�Ԫ�}[ PD<�&���U�\���<���9$�M��%���*�M+ػ��4A�Px=��$	&3�T�o���q{9m���@G"��x�0}�_�R�WK+|��OK"�١ߛ�1Q��X>��l��@��h^ȵ��	��'�Jh�I��^���=*��w
�yH�㛄����2��!��?���s�f>u�)�߯����f��
=�tC��`�Gi�>�����'_���\sᤍ�-�	pkMIC=P�y݊I�IK��j˸��U�&a��W�֟�
$���{&���@�NsV��W���tHBkn�h��ʘ�⇺��A�W�!P�
)�l��y���f�Dא����}����{�`k���-vX��O�CA��
K�Ї�v�ķd¢��7�� �~�5�@��x��T���!ט��ȏp�M�I�F���0�F"���G4շI�$lդ��j�<�U�#4�V3���6����/܏�yU�Sl�l
ܵ���|9iK�fZ�NF3���T7���'��}Y���L �'Mq}`��UA ط�܉�J��ɮ����	�]bk�E���M$Z�rr��%; �	�L���N!������Y���X�l�˜"^���I<��w
];�_�/ٴ���O��\ar�Z�:ɗE1/h�_<I���ٱO���AHBq������y��M)�w;�L���%���\���sm &�&Q��ؚ0�T�+�u��ywgٶ��u
��!��U:��Δ#�Y�me!E�F��0h�/�o#��\e�g���A��T��s�X��O�Y�A F����#���`�����?r2���b�w�\{�ں��n`!��S�d�W���c:�e~��LK~n��4�9:Ł����i�#��]C�|��hG�±ߌ�ΦdKL�6��W��j�3&(b ���l�pGRA��2�a孶~�HN"֒�����iH�*�WOWwyA3ܫ��2D�R�:�/sS�u��	+�ÙG0�	�uotc��.����p"�_&��i��/6j^ʉ�ΘU�-<5{o�=2��-��h<����L�z��|��e�Ws�X��R1k��^[Fjp�����V�zzj�3�"҈`�*~C%O�}�/i9JꂊB���d��F�����]�%_"e 7��Ԍc���Ɩ�� ?�TQE�qy�]u[¼��j�<�x� �Y����8���E��3�ѳ��1��w)n�Q�� ���Fu]��a�[#���9X�اQ��R_�Ʋ+�X�;ucw��o^p9�+J���b��'ظ��x|a��]>;:�:h	S��hi�y
���|%�6%
�IE���j�B�C
.�b��[��ۗh�E~4��J��	b�C�/��5E�����wwQ0�f�|n$������8�����;.Ą�a�[�y�������	cR,�L���2ܺK�>�ׯ�>Q����a�$:���S���ϾpHH��k*�٧�8��� ��.|�~O��r��AE&��I��iį� ����^KH%��w�0F]A���2�]���<r�R���'6;�C������QHW��J�/5�������M�SS聣��n�����N�˹S���fy��nv"�D�_��@o}W��$^C����<�(��z�{�p���!�'2�#�~�4 2��[�Q F'�w���J��q�TjK����/����RXlxVHYEB    9620     d70��~xY�K���u��>�!�xkC���*�7��2*W�lb�ڌl՚�D�'_<m��7MP-wXF�1��!�:�E�qM��_87�st����F���NعޓBr-�H7����q�;W{ s�N�X���N9R����;���q-�Ԭ)̃y#hD��C�03�������MT���+��
�z|�lr9�a֋{tΈ�v<�A�;"��\탯�L���OxUpeNkj�5bYh�d~K�d�~i­�uf�lq8�K�"�b wH��F\��3b��s��t�5�DwQ4J{o�E"�������l垸��7�ʔ9/n��lc��o��o��`�US"OI��p�;.��hP9�9���Au$��-��.�A_$� ��!��O�\�H��ƺ�u��
p�U�-o�"p�*�K}���>�B�([\v�S)��ա��`�PG�9�]mL�K�m��g�ee��ɪ��g�U���̃�)g�k�\
��6	�v&���'ޜ�}�Z�'M�_��w��8[80�a7���a��E���Q�3!�o�4��*�c��o��)�y��1z��B;0���R��8���zd%�&������<�ʍ4]��1��:�U��uP�Ȼn Ֆ��2�94 C�䏷LO��\����x�S���c�@��F�J~R>���&:=�'�YԅȒ��9�����J���<kHL6Ĵi�ey��#_��jm��CB��Zc:"�\zv��=˱Ǧ,ȼV��i��g��S�Y-w�L)�L1X�I�f���6��K���f�bq�W������b{�u`�!�����kJ$� ��K���3�M��+i�S:d�,�p��ӥy�I����z蒂�r�{=?�~hDe9l��B�;\�=7�˭�y	.��5��L����Q�~1��1�;
�}�a����-%F���`k�j��AX���$v��Q�ߏ��A���(�l��Z�-�\�{�
���ba5b�7�W�=2qm[�����Rc���zP ����ned���E��n�!��N:n�9�D�$6,��i�ǝa��S���79���e��7l�~��ـ
.�������P�����M��G��Ւ�����b�IF�6y��5Չwz�Θ���j���\h��\��	0j(�h%X��dq��Ⱦ������,�l�፪�S�\���.Ř��)$�)���~����K~6#�?Ď��>H{�9��G]ծ�FB��VE���\RwV��p�:|uD���Glt(�l#���ߐ����	ٷ[������\�RH�q��좲*b�Q�a\�Ҩ+�'Aa��W�:f-�n��	]�뫾
j��hN�q�N)�ֱC�K]��Â�^օ0�B&?/r���߈��r8�ƍl8ҥ�dx�s)�4�̼3
���\�����f� �� ·m��s������[%���=,_j�z���c��X�N�|,�b�
��^��Ӵ����8�ޏW��na �A�X�+yC�O�rĘ�;��HZn-L�V�vx i~gq��3`�	�Z0Z�������{�^�VXX��]G�a�̞i�6p9h��*i�	r�χ_(t�'.�ћ�K|�qe������䶖�+�����q%��d'ᦑ������6eb��rx7"] 
@ۑ�|�����i�3�(��� ���Rd�[�Gd���'YS؆h�:'��.-�x��p��zV�S���>��Q:�<�ދ�	%�o=Z_�[l�u"��t[؋�Ks����ڋ��y��Iaz&x��v����J"q}Mc��3S�L�Y�A��g������02�,�<��G*{w�C��6���bN�<��2����|j�e��ꁯ6#$���_��ـ7��̄��r���T=P�'��'C�����{/
�ŷ���jp�����s?�~E$y2��Y��a���������� CC�*�9�����]}<��0���3��z\�5��_��r�1�%��=��Yd�PW>��t^�iT�e�0��ߞa%f:Xt�"J�6Жg�����f�
n�Z_4�-> �-���w�z��0o��xgd�@8�W����:h�:k������@��ڛڝ���C�ă!Q���5��L�y�7�V��b��/��s0�|@G!��ͥ�
oH�Z�f���T�<̏�{��T��^�,�x�j�4��0���.�7?~D�Y~�l(�h?K�`
m�Q�ʵ��v�^��雂)�ӓ"_����P�����&n��7e�|M[�=�ee�܏s������:��@�ʟ�@@�n"�T�,s���ap�g�����7?��(�-y?�V���F�rM6����FLUL�w�<w�.Bo����vLی%��\��a��J��_�?e����rtvF�𺭯��z� �����B��YN�#d$���-!�A�)�̪�ub��|f\�'U��A���$t�N�ő&��9v�đ�DQ; �v60��(�����>m��:D�~!1t�XX��y:�$kSg��+3��;��#lr�w�nɫ|@B]��%�S7����~ Ѕ!��w�4�`����yo���Ĭ��0T_��t:�����cU�gs����Ir/(�.����o�,$��zR4��p���oܕE8�:����}m����EJ�7z�ͩ,<VJ>^�Yޠ�|<V�W�Z(�rH#B��zz�o��W6f�6;v�� ��V&p��Wx!ة���j�=S��=z�]����t��P�e��8��>fS����ҳ�=%�>��>L� �@�2R��so��|�tOlb�o��BR��҆lS)Y���*�(�Ѳ>��D�\�sm���7QL�z4#6(��ɫo�~��L�OY,0�T��@4������E��3~������'No=8�����#�>_h�qY!�Ϳ�}!������1�%����̎$�3)��$�|\��~*�XrJ��3͟��4���{��f�����&
���ղ>wJ���RA6�4|�.Op�}س��Z���W�U���  �ƔyJ�
���b�Z�WY���I�o	f��gM%��JG�gv�v�DtE�/z4�"��p�a�O��A|�%�5'e�!��c���T�n2h�7�C�R�`�Q�;S��]��9�N��}��.�:&�mU����T�)"]1(�3�E>`���$I�ʱ���U"��P�K�)*�1���E��'v����~=A�]��"��Nj����&d��t�JѫY�#����4��m1ZN%��✭��Z����*zeЗ��&�����D�`��d�I���VYj�BRť�� �L�l�	fc�LOK&ئ�y�Y� 4[�2�{H�ca��K: 
7�<�QO�ñ�ۑ�����6�H�RQ���@G���88?5��>