XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����)��yO~�qǀ�>�~ڦB����4�����^x��G�pY`��qJts�]�����><�/��Q������i��пd,�W���K`heAID0��9�r������'�~�Y.Ҽ) T��Ĭ6v�P�d9�k$�G��R �鬼<)~7·S�� JE~&A"��2,m��q�k8�d0���G�������az�C��L�#(�x�C�EtvA��d�,� E�7l��|�G��!��LWH�ǈǆؿ2�$��ꄛ/�]ˈ���صV���$g��Y���� JӴ�f�n1��ů�$Ur����_7�3�_��Ȟf�T�R��i�����x7�T�J��<�]�������?%]��g����q�\� ���K���;�Ფ����@F����|��퉣���v~��z��X?�@*q��y��U~X+��,� ���ko�4�D5$��Z���C�������O�׿O��:ԍz6�*���N�V�H�ި�6��/�:�w��M{�%4�
�s�M��ހ8Qm
{�a���G�$`+�0������P�B��Ly%d�9*��1N�o��GفZ[8M���fy>frH\�H�\+
��_�|.�U�����)��`!��? ]���V�}� )��� a���3~��Í�Gb^�3��W�U��WI��e#P�ž����b� �VU$�|��{>���M��� 4
��g�?N��F(���۩��:��x=G������Z��~XlxVHYEB    b8a6    1ac0���E�J}Z`>�~��:���AY81������j�ѥ��0ϥ�����.fkI檚PlfLC�p+ߚ�Y*á�B�h�=i854��ְ������o���8X��o5�lk��Ԙ�):�3yH�֝�&��ܒW���!�a죫=_9�| ϱ?��B��{'��l�"�h�cv�&��Г���`�V>��ȋYi�	���;qP�I�DR�Q�\�P�L�.}C�2���ekpռ��A-�n�!�x�=��Z#�Ga���6]ҬU����)�?mϴ��=^���1P�H_)�A&\\Kgue��Ӧ��7��םM:�8ld\ǵ��WWl��9g"����J/�$�zE�$q�$��]Z��T�&R�$��J/8���I"+!�\*k[^k�*�d��!�p�M�DU�����g�����!��[���˙� g�� N�V&�6J�������Ѡ����8�nP?wApp<؛�;�(�;��1m�����v��4j����%��L���ڢ�;�����e�;a�%_'�60c�M�6���9�P�_�<T���ڡ��ֱzE��%K�Rՠ������\�ꜳ.(~��1�fw����|���)Ae-N�^�+!=+�������53��#��1ݍQ�&2����l�zN�ÿ�m^!Ʉ$�=�W� �l7R.	�K�vbpIc��M�%���������|�Z&��$��f�>J��W<�=s�^'�rb��e��ͧ�!�4�*${�����}�^Q�Z �WETw�y��/�����g�}Y�.5��G�,<)�a4�� �/��a���	t;�{�ޘo�a�آ���8#�9��2��k��G��3�IUM~�����=�����jQ~ �Q�t�;=�h~����zw��<{f���Xo�iPO�#�!��&�s��m���͔O��OU�e>��Cl�XBZ�^�JMq"/~ Us�<!,ƓK�Bg"/G���͏�i������k�4>|;�k1�����u�@H�XׇW�G����)+��V��0��^m<���S?��!Y�X�q{Ѕ@�R�@�kv~����^���#�2��pF��0�;Y�An�}�հ)v�C$!�1�,��7ԝ���tf��陚/�}�`�m��*�L�VN��2��?x�M�O�1~�%y5�/]i�����%��˪�,�mi�9����*'�1���?�R%�=�q;��M��^�����'�އ����U޴��s,_��^ �e2r��*�{�1
1�r;�;	���-��hZ��ĭ�Q���#A�Dp&9��t�B�`]�OF��ʞ��W��H*���MQNw��4v�'e����a�G1,�I��$�)���W���!H��
��j��kێ��a�fe}���Ηr���,-��Y�+a���K��M�<���7�f�tw����f��ĩf�t��Oxe`\|��E�:_���@'��3���B�0�$am��D��1]B���|/�sV
����&ۜ"2�9�zy�T�-sÕ�k�#> ���Z����d�+���4��������2&��>�^����e~ �O�x�ɑ|����f�hˮY0:��EΞᛡ�Ƣv���-�綏�(%��dgm>����㰄	��m�1?b��A������I�4����1J����q�D�;'�f��M�(�:�5#������F�r�f{-W�1�Q�����m�� Ի���"�x��W7�������6S�xg�Oqy%(���$O�l
͖��wDy���= st@S�%�ӥ���}��}�0�BXل���p]z���	EJ��״&�_���M4�����I�?R�f���]�W��G��=Ȉ���XT��}�N�Ud�.���L���k���PV��-�(�"�?���Bā�
�%.���w�/ <��{,���=�/6�^�7�촩Qa�~�6��o��^��vE�҉��� �j)��gF��ۄ�h��W���"��&�`#d'�V�b9j��ߞ	6�;�1�9J����,���@.��m	8w�Y�84_;iZ������.W=B�=x0r�h=��;�S��cԍ�������:��Gg���γV�*�S�ui'�@f_�r���1\�\�"�O�A���S�����د(�Ɋs�>��77r�q�2��u�+���;��ܑ�LDQN��v�� �ds�������DZ� �����lt@���)B�*R����tCi�_�Goќ��	`�z����`�m��⬗��/���10���	��QS8���b�|��:��Ac�jù����'�2�g�%X�����=��t8��I{n1�N	W�´�)}��^��F���t���	[*��l҂#�J�	�e_��\�ƥ��z��l�.m���G���AP��|lf{��Ud�����l�u��3��s�Cf�8mc���#�	��¼֕+�HC�	�J�m4\��z˗T�}�<��a @��o�okSp�/ Su���m�a�fH��髅0��Ϳ��ς�A��)�I�s㝢Q��U�Y���deJ�9������9�rػ���?�tq%9wg��>�)�$��i�����?�h�7�v�dґ[��9�� 4����ɜU�oq��=Q����Zn��QR�c01��'�	۽ !���������r�vެ];L�ZK G,8T���4��io���X�?^'�-�{�� ��K�޳8��o'�a������HA��-���a��RW��������d&8�ٗ!��;s���UU�O�ژd+?�����+��s�@6f�3����S��i5�R���=�؆0�FD�{E�	�,��u��N(����ǣ� �h�0%��S&�3����e^�ד��WxFD�
gX_�<7��j�6q]*�1�Y�5g�WU�j�\T�Q{Xh�g&��9?�^-q�wI�x�):��vr��+'/v~��A?����@���"��0����wt��=&���7����͇�@Q��B+FBOf��s4{k4��������ku�+r����[JI���0#�Ȩr^I��Bw$�/�~��9��=�wՠ������'�t�n��j�^�4����%��#���2˷ 12�d�4Vn��S5Tf�\A�35q�6�E�|H��ؐKJQOi�J����zꉿ̻j��KؠnT3�}��$3�L�'��qg�"���jLR��"ϋ$����<$i$����?�GN/6�X�m��w5�j4T����5��`ڮ����Lk�60	ҷAM�xH�����P.�[2�|�I��z�V�PX�!g�_��/	�f���
��*��I+�̒%�>��z֫
�  � �1���{՞XG�6Jح������`�K5�z�63����`����p>h�Eӌm�� ���;�,3O>��n# �8|�"C�n�?r�'
��A��4)��<�������m���Vy����r"�g��9V�r[�q�����)[�����������Γ�v*� ,M�׃��u8Z��|=�,�S�}Qҧ��e�#�[`q���y����v^������/8�P�hY�V�V	kq���b���߮�;�//�'l���pzɾ�������E�R��a�-�Ĕ�*3+���ⵎ�a���O+���Nl��V�&�����L�������4ȣ{.o�D�+0�k4#-�Lu��3�F|��Dr)���M�`�����^U'6�m!Z��cD�{���?�r?x�=��i�u�j�8gEȟ݋^�Խ8}Ɩt�_QHG����Y��?�R�M�p0~��l�P\�|>��V�9ďض��� D�x� �ЄJq�)�u[u(�d�|���KN�?�6+�pk������~��b1���_�e�:,d�(;��S�� @��I��@fjH��v�|��u�G�O��R�����/�	�������Z�P�%��K����{Ӻ	�t��~�Lg?�Ղ�5��	��\��	����5�I�Ho�=�v�2�I#B"�j_L��}���s�l������E�NPϺ�L~�������������&�7�))S�l.j�,�[�C_�>���g��[�Uu�eז��(=�)��_�)�fS�j���j#ze��/_�>��|WOj�X��/��ŁH�Ykɿ`��l��v�J�)��@ �Mk	���e�*hK�.�o~?�ԪPq�v�ԞR`1�"~y)�c�Q�aH��<���:����Tk�eL�T���P�&���oc��@��jD�,x
/�Ԫ첣��3�1r�e������/* ����fT�N��ܿ�O����c`�ŉg�.>+C�9�$���i�@�wז�4-��o�����V�����ʂY�jE������|0� u?�'�$E��������c�����ŷ�x����F61Κ64z�Ve x)�A��m���[�`<�@-nM���O����we�( ?�2w1㫥�"��=WNlI���G�&�ɐ\�;j���Hh����R��EK�L�R���:���c�q�����*�l���tS��%j�V��e��x�c6�����FP�nɴ��
����$@�(O�%
/wni���|��2V�y-u0��?qE΋��8��Q�VXB���3��L�����}��$ώ9�G���*�
 b��͆P�N��4{1��I��{���L.\�2�o��������"��+�^����t7Zb:h&bt�x����/t#TCF77��S��+���S�7�u�Q��+>���.��@�N�f�!x����#qt�2�E�o�ȶb�������D�� �n�Y����UJ��A�&���I�Q�c��H�zB!�*6�c�g�&q&|��Q��|�M}��~�MC�+��Ĉ����a��'��H���%���Yhú�H�hp�+�w��ORrUz\�|��s�K��:sXGC�9V�7e�S�K:�&iF�"ӊ�9���֏�� � �u� �~#]�X ]�48�1� ��aš�ȆA��X��$H0S�QZ���R m���75���WE��=�jnI]-��Y�j�YR��N����<��n���N�� �
'K��g�����k�@J+m}^�"��3�X�dkPf0+?�=ܭ�ߩm7��Ά@��KԎC����vV�)0���,��l�8�ƽI�1y�lR��	h6��6d���ɻJ��>�s��&l�|*{�^@䤭��`�I݃cvU6�μ����M�%�ݟ�#�W:	4E�0�ƯYP;?����* x L�ӟ�_���ocUu���X���:�R����U����%�nә��=��g1�In��1�O\�f�������4Y�HW�o�,�\LΘ�;J,T`��]���)�	��z��u<g���@���P�m�uղzd�T�Δ�\m�l��C��Ǟ�D�������P�*@#�]`�U,��);�e�٬��r��m�.���t\�Y��u���F���5�Bsf?��f�'5u�A���zOڮ�<��Pxֿ�l�'؟�IN�O�R�5�@uHS���CK�� 7�"IolWW�]��x�i�GhvT��ϰ8�奋��.�Z=�3s	p���&�6u�_\����r��-uC�Ҩ�>#%J4�q���^	4�1�֟�ʗU����i���ccbt
$�!�dc��䇷=eݧI�!�2NM�f�u�M���b4^��+9��]'ե�	߽�틺��c�«5�E�E�2��y>̺ԁ����b�#0Ï`��a�����#���>������G��_㚤T3n������(�F�ej��:n-�ȃ5��/F��II�EZ2oȶ�~���ࢱ�6^wl	:*\���]�ٙ
E:{͜��Y�R�]\* $#_��S���v}�ݘ�(
�v\�Q�v�dFZvy(ro2Xz�xٟ�7�*t�c�D���< ������w���(-��#y�I��eH��B�/�g���h!��p�y3{�!z��
5/J��)[�v�l��j�2�U�4�,�t��$>IY�{R�������aS8�t��<�)��M�`Y��6��R�>t�ǥ�pĄE[�{�bR�GG:��`6h�*��x��')�K�F�9�p�������Za�B��ȚG]S	������`���)i#Z��o��|����4t�xR8^���T^[ڇi,�~/�_�e�����)��]�P65��/k��(6���Y�f�D6�cJ�%�W�lþ����3���ȃl�Rio����������A� ���bZ����1T��(�N�&K�l�//d��"p*T�3�>���L�Ƶ�L°*^�v�B�HTgB�W�>ɔ���z��E�=���(~n����!
S�a�'�%�`^�x iC���-Np�h�Ŏ�,&Ӵ��nJGǯm4�u� إ��/6Mf�x�<m֢�SPif~ْ���
��~g�`)����f²&��(F6��I����w#�-m�u�U�����fG*hϭ���eē/.�_��X�詻Zj�.Iؗ
�֞�v܊�����`0��%j��
ژ�r����},��Ǘ��W"@Z�1]
DCmi�Đ�k�9e�cor4�c<PEC�&(Nk��'?�E���+�Y�3e�� a��2��q)8��3��������Jf͛so	�]�N_�K�2��s��N��И:���GԿ����k^��ȑ.����>�E|���icp�w���G<�������+�*0�b@B
�%C\�X�����:8�O�`:�@