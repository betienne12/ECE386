XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������4����)����7�������iڞZG'�YVe�Y_DyT}4����(�upu��6�\�N{�%q3<�c���pal�cF�����q��<�_���=jΒ��S�#��~il�wq���_}�P�s1��&��y�'(m^�w[�:]�5Dl�0�c��`\0�cw^�R�"�y)&��K*����&����>��Q��H{T?#]�e�ڶ&�`?@J/Nv�ފe�0���ƀ�	����ؘ$R�������p�"Ř�v��z���#���4����7��ꝉ�d%�;GO�ʂ��)��Q�{�܏02 ��\��s,��r�J*,'����FW���]a���}/5�l�*�����6����1eSޮN����f�<��ߋ�����G�\�/�8��y=Lb���v���^�s_����ީ �,�<鸓\���Bf�����Ѝ�3/���+`��hq��$��p�ː���(~�%9�8�g��}���������*�(�u
P"��v���-p�Sz׭7]6z��Q٣�f�u���f��%FY�?��жJ߲}Q�����^������2�{.����7���5��?� 8�*sMw=���؋ G&�N��<΢����*�����WO+�駡����BD6̀(r�4��iw>�ljo��
ze}=��kvu,�.��Ub]���6`OC���]w^�U��5��@��V��a�rN�0�/���Mg(6$��Y*��0N`u�W�NfXlxVHYEB    fa00    2950��d���L�U%0U���e'�yFnI؎����C�j����L��9�����4ģ�*�ԽnHL
:�|�����t�S5{j�{�t�g+�dU�Q�;s�c������p���J��nc��b�EH��cmZ�ZeOn��	��7%Lф�U�����n����ۍk�>�'�7�8*�s�����I0��c���q����,�?�4�����h� )�*>�]HZWI�,b�h� �GGz�u�E#�&�T���yI5����� ��K~�]�|f>�����JU��0_K�&���]���$8�u<O5�]A$�T��'���¢�B����P��uEuI�i�Ɣ��f�$�+��kN��}L�0j��֭W�D���h|�	�>�&�x��N�z��4�'y��t���g�0�TC�.��O�i�@T����#Q�3�"��7�!0�,��\� ��?�r�ײ��S�n]�����,^J�p��ȹ�������m�.�x�,�S�ʺ/E����F����<��Rm�OJ��'a��M�No�ZTI
T=�e>`,�_M�@�j�)���ë��j��
	9oZ{�K���r0s��s!a�v�T=����mZ�T��UZ�U�eRj0�����x�_؋߶?�~��gmySȦހFD�����-9��k(�����i�_�ӈ�_^�_�(%k���=�uc:|~�Ey�����K^�u	��@�cދ�!x�7rު����з>�kbx�������$K�e�'JC��5�)ǧN~�$qIq�.��:P�&�)���|!��ӌ��{���y��W���q��a.=`����X�z	 ���VP4��$�p�=:Fj&�c�q�7N��
0����~�ؤ&.�?ݘ5�[%�1#�� K���ҟf�a:)�P�O�$��)��n|:ۢFƻ]���mx������V|����y�K-�O%LXRa�Y���BT��Ѫ@���s*����R}RX�_w��(�,u�]ך[~ ��#��s��گ�Slpu��B�(��pѼ��,�/g��j퍝E (��(������W�'"N��Z�w�����*svS��kb�S���VR��8�b�/�/�|��E�Ԫ�G42��Hr����gsr��}���-�JYAW�De��'-e9����(F�j���`𭕨5}Qİ�@W�C_b��?��Z$g�q˵��?l��#�6!rd_�Qs�]�Qj��0��w� ��]�]s�- ���F������9�-�n���,��u�C���y��oC���n�1��(_����io��Q�Y�"ud�aH�_���:�S�-VWN�bL��dD�?Tt�vۧa��A������G�G�w���� � BN�uZ^��Q3��UH��W����&�䜔8���zHSb1 uF�<f� �Jo�bs��$��KtN�,���0�������h�_*]Z��]����hD��� �m<����[\0ö�,��BP��Ҧe>��Y���j�g�Hjf�{��N� [CԢ��{�9�>1^$�F�8�-?*zp R�S]C;��7Ɏ6�ҕ��|%uOǼ�7���8&90��U;a��#�,�Ek	��W�=P��v�(3����vO�hma��2���]���o�?�A�w�.�'�V��v	6��Q2��2�J0Y�:�̩��G.���/O��2LD��y�u��� �8S	�l�5�\4�a����.�f}X^�\�w�ң�&B�2�$�MC~h��^�G�"ݲ9��v�cִ4�E�rGc	uOB�CytsJ�td�OAn��f�|k��ڃ���4Z԰��,��=&��b� ��s�@}��|~�?P�Ír���
N�*KV�8�
�v���5�'�a�r�~V��Q�̩&rޓ��6�7�G�13g���.��׿T��G(R��������$�$4;�&�wy�dw{����p�U�$�/p��2�`��c����dtM.1�����������골/M�9�/F�ת��d��oH�z=�p���]+AM�~�z��]�f�f��P�W"7��E�xD�_bѫ;N�q�d��?�W{�l��f�7�4,ɺ3�k���bO���*�H{��P`�y��y��m���|�^�#�z� �U�2D����@�!����7����9:�F_�_{�P򽚵Z?#+���i��c�[��N�����YX�(�a~ۏ�]����M�^[�)�v��v���
l��{@a�������&Ǝ�Ջ������l�Ol����<�@���3�g�sn���������ض�?T�ۓ���Q���6k���h��Q�J��=I#Ae��#bv��/�V����Č�Y ��ݸ��2���;$��󶬦�4��Ko����:LP9a�\��H�n!��y���.��r���o��9G�a��sY�����_=��8����x��v#��k*�E��>++�wO~ؒy��Pd�K��.���I��_�Y�u��b���� w=d)!���]uq�g�!�C���$g]O�bo�Z��蓨��N�f����5ݦlqz�C[��g7�~����=�X�@d�a{��JkQL[TT��_�J� 
��P%`X��߸�\>�Ve����ڰ�.�+KM�	у�Eͭ� �Xi!����'V�L�oG��ՉMR���v�F�<�9g��7�Hg�B������ �(3�'f~;�gu���]��s�����߬�:����Xl(�Y#m2�Ω�g.���������H�o��b��%%�k�6.�y�5lv�e�����yk�^��L��.x�}�zE�v�r������G.���@��f����^J�����������,�%�Mv�rg-�Ռ��ϸt�|�3v
-@}���Ϣx���A��bG�=�sY��c,���'ӎ�)hh\A�?�
��M9]����UNr��F��e�d�b��� �F�O���4��}I#Y�Sp��||D~��?��/�)4y��N�� "wK����r�{B#Y��Z<9�0���j���������vL'�?�E&��?���b�������$���7�5�'q:Ӕ_Ĥ��Od���VW�S�"9/�w	��κ.���vi��/�W�سTz��Hj}�e�Jrֵ2�X��G��u��r�}ְ��4��ZdLrG�"T�U)� �ٝf���Z]4؉n��F(X{*K��8)s�,�*����L_��x1\{�l��05��\����#p˾��;Ux�~�Q���5h�[Z��Oؐ��x>��.2��c��(:�A�r�9l^���A��}N����THo"��y��"�4�sf�3�$Ay(gS�����{��q�1A�@Ĥ�a��˕�m�pC�+z�اS����I�b���P?xo �z�U5o�=# Y�^�>�73�+�"�
�j��v�v���{����m�G�t�z��sQ8�{�.��`§�V6V%�;Dl֓���Bb�c�y�����-x'GY��XK�1,��IWa`���.�ς7�~꿂�)�7U@��,;��<ѭ�mw~��)3�>ڐڳf�?fo
?�WP�nQ�cq��}��2RS��N���`��R2�!)E�""0'�٢T��q��~n����	�ȑp_��;���i?*�OEx��;6���5�*b�C���*����)�e'��M��֑�z�,�B:�� {��N�'�A����ŭC������/lG�o����*;���t�V?��|Z.�y�W�B���F���T��3�Y��v��n�#L�J-0�6����F��7��a��}EeBj+�H\��E6���rye(K�E�ӗh����wlw�<����.)�+�tm�+ZO�9h��1������;V��,L��*�V���μ·M�͡�,��k�u,�*�Š;�.i�cR�?�J��淤��3h�%r��� �^��,�?h���#4H}w^F��0����@��_ 7	���N�B꘿93A.��`Q�A�/���g��DAmۿ+8����<�Wu �B?�*e\1�3]��
E�w��	+��p�rY38a��T��Җ��Cὅ���;?D�f�#��*��H<��5����6�C����v��7�i��̬+P��Q���a	O����� ��Ő�:�~�I��K1G"�T�	fSq5�f߀�\{�.�c��Z"��@�������}oP7J`#��`��2]Q��,�o
���s
\-l�JE[9d�r;���ʞ��k��bD8a�ɞv���~Ķ| =ƿ0 $��{�a>�"����:h� lɘ�P��c�d���z�Hp,�L�K
��Q&Q�f��?���<=��|���M��0�z���B�$KA��$���cs��>����#}��h�hP��۔Z�� K`k����,"����!�N����GnB���ʲ�\bf�5��(�C��ѱ��d�W`>���� (�~��wQ/F��T��ֶ[�dso"�� '�#>�k��?�0eC�w�����Y� �w?�]����8v��]�Az�q/I����Y3�W��Ηo:,�b�:��d�>)-ڼ�e+�} #h|/٢�$�3V�M�X��Vy5�.��[�?[D��щ#+�����4��k��n埌І��^q5��)����~���'c�.C�XR��H�C�aI�,���R��� �:�[�:��(���,8�0�{��}e�wZ���M�W�p�k��/��/45�e�;I1�nM`�`]1
x�m�!�C�/���Vh����!����1K[h�֥���f���-@e��믿�p��`@(� ̞����S��.�?��%V��O���?�xuS6$��vo����	�?�����|N� �=$�����M����ܠJ���B�l��t�Rq��Gk<����_�\XQ�.���K�U]!���gO��xԳZ��xy�l�xtEG��=��,�w^��"�. :�����p���䩇X��ap�ǶyA����:S�VNK,3Ґ%=B���&z=P2��a{)�yɧ7�x���_�N"E�����'�8���5E�`%rG}[y����J�G=�����٤0-�eư~5��Q��rN���~~H�ER,G=m�%5�����`���3��N��� i��jkn5�-7l��6��#S�tN��2f�q���w�L� ��؈$ƒMˎ�Oҗv]��L��:�!WE�BJoW����{�p	��ċ]�	��/���tq�?�Â�3��Y<daA�{͊K�0��� #��?�T;sѽ&.����D!~,��&�{�c��@�*I�$���~���cu���-j�v_�<$��2�X��V�M���Q��<ş(�糧�~���Y�7�y9�{�Ek�e���Z���]V{Kf:���+m���G�W8���t��e��ǰ���l�3�J�{�� ��P����K��X�:�3��&�k��b7r}������O"�H�q��!��r�Y�@5#���ʶ	�u�y	woG����q��(�?�����3i�O��U�j�&�+���0$@�KJV��0G^�����5c$��k*����,~��毥zf(��(0!:��Q5��_}O���߅pă�+f�e�*"Y0�&�}����)����	X]��z�C	�Y�0>U�߳$B,����k�	����-G����޴�Jכ<V��c|�ؤd-}�����'n���P�!Xx�|7Q���'C�a�:��g�|L(K#m��j�='a��,s�hh�OV�a~�.�q,ۍbxM�
y�Ӧ'�P`��]��9�H5���M�x�f�4�A�p$3!<�J�3���_�5A0g�G ���c֛�V�E�e�+��}7��_��L�|��+��x��n:'�<y�!v�H;�����/��_^\���&��&R�\����Vj��b��|�`�k�z"��Y��̰6�{�HG��#,��K��8HitX������]}<0����\��n����L�i�eL�r�x�؏e��.3��$�ƌ�:�&bS�^� ~��W��*v4k����[�l6\L:��Î�Ql�g�?���8{��������Z�=Y��SP��l_�����f������R���2�J.,��N�m�L��=NW��Qj)F�S-��x��g�y�<ֻ]���z�b�/^�9��좘����e�3%e^�^���jO�)Xʺ�L��q,�7r��P-�����-����뭦���e��]�Ǣ5,����� }����koU���O�	k]��VqĖ�q"c����b��V�L5���}�T���B'|.2:��$yU%��W�Z>�'�*��a:sk��0b������Z3|��<���B�LSW�'�
p�������uqZnm����`kA"�d{`$�H�Y��9	N�/ھ5ȍB%�N�qэ�h2"����5�Z(�6tKn��e��c�Y�:m�xj�P���� C}*���*�Q
GskL)���D0۲#��Q�#��uHe2�ǐ�l3'׃��0O:�����K�A��N�8�F帲�0�9���^�h�����2���Gao�ʩ����е~~�Wc��D� ����(�\���`����^�r;^`�ofe��0/�a˥�a�s�u!#�k��d-{;��۷Ns�j�S�!nnv<�'gp66n�[����[��P�ZE\L�at��T�~#
�ptz:XY�E�����w؋�f����O�un&�}��eU�p�7�8"�W4Z�1�-
FP�v�[�+m�������aF��k.�3�S����ii�����;b.�� /'����}NK��XI����Fk�bO����"ޮ�&p����r*�#(�H�%Ď��3�����?-�6:��C(�qg}_l���V�K7����"�����KPe<�q�^F�ܥ
���4�]8&0��I����K@����r ��Z�T!KB*�j3U�zO��/C��G��3���r��ѝ\��}���Ai�%�ܪw��p�[��;�B	�<�nHh��p\Fhy;�[\�3� ��z�l\7��?�Y�ln<!b��Cg5C�m"�g5��%�&U;��6�}3�ŪW��V���PB,iP������� E���aH};�J��ܶ�<9�bk�f����&,���G�m�[Nn���Y���b�*��6�財�F����F�j�����2R�l���Ol\�4��̽H�72���@���������[,��#���\n��J�����5:2�{��=h,��~[�"�E�C;�!b���Y������d�tn띬н�·�,F&LB���Rz��0��g�w	�o ����}�ܳb[�>PiX�Q�J-�湜�b�c)+�Ճi���~��:c"	���}�W&'�
 �Q*��c�--�yzG����rq�-�ǭ��-ʶ���3ܬj��L_�[�\�����X.6�{x̗�6כBH�Q��^�N��f����IL�ic��;�%M��`��R&��JR�Ć�����G%A�vU�+��{s.�ϑ
�)������/����	�>
Y�hd+�SЫ�4��%)�=�rx����J�Z��ؚ�{c§�5|07�� o�?{���h@u�Y���$� |�MɒY
����X=r6��4���	����4k16S��k��)}f7���.�����C��&���}nm\��
��qb�U��q�&gc�
x�P��U���b��Za7j�!�a�ߴY>�;!��i6(d����H�8�S*�s�T��~��EGu��u]�M|��;�^+K�w7�d�����@;�[M��P�8k�B]4�@�f�G���e$�b�g��my8�l�y�l;�(h*���W#�0��G��F�F=>����׼�����ጨ��FRp��r��76�����Ej�����
��{0h
�Ցi��8���{r$x��C�V�[h0XɾS�;.���<I����o�y�i{~�F}ʜ�b-�I����+��������}��?���,Żz�T�3��|�&��|��*�-JsS������� �8 �Ȃ�_�*&��|�ڭ����ΠlV�e�B���F_:`~�:�����v���ڟ�M��1D��Sqa6��������U�8;%�h�~9<�^evsY�Kפv�W0,���X ��^�+�#6�v�	K7��ænK6�T�Z�.�����?�i��'1!L{����{�*te��H����V�|q~���e���1]���!I�>d0�+V�h��(~����ĵEǦ~h��3l���C˭�� (�I!#�M|%�x�#6֒���V�M����V��frâ��.w~\���?�3���M��/|����V:�����j1n�!��wDn�� 9��x+R��)�c�qE��X��0�L1W�K&�9�bG(f[!7��O:If�D)�5���7^G4J�,���a����\���{:H�`�w[L�K�UD9'S�;�$ލZ����`��4�>�B鮸^�ptB:�˧��	T�ߣ	�R�������Ij������@������;ܺ�j���8j�x��lq��Na8d���5�T����C3�˷�!��pi:��ÀGu���dnC��a�	 ��D��!�[<�� mDG��i$�ՙ��*�1�B�f��Ͳfհ9��̶�Io=�][]��;k�^F�ʑ�Py���7G)��?�TŘ�x�L����h�2f7@�GW8�8�]�}�^PzpH��0�	6��������������&�\As��)A�11�Y�O��q�����PATJޟvfמU�`J���<�rr�4ɲS+,��(�ѴHpO37
�SC#w��+%+���d��+</��ka#��~�����*,�Y:�7jm�po�HCj���a:��'3�I"�-U��|=�+��D�����e�1m����ePupu�ׯ�@�����;F�Y2c�`�*�,��P�A/�Y��r�����f�G@�����1Q�q86��I���fᴮ;�]��h��u�3��-e�R��VIK���DvCt1�TT�ϙ�}n��\A�]d��&
i�k���灌���˧���Y�z!�G����]ӑ�i���3�|^v��&Y���</�J���ʠ����g�f�Q:^k��
��.�����
d4���
,�L�K& ��eJ~�����F��������5Bz=�o��CJ����!��S�^��4n��#�(+� ��Q� �ה2��U��a�Td�(���<盿FD��.+;��\����K�a�����������4>0��,��zM�mEUC��ߜ�L��(�2��[�P-�E�n�Ŝ&5�5�p䲨0xs!��quQF�[��·��8V�8m�Z�� x}�_�;��eC<�~���,�Dd7���_B|��j} *�ܕ��/�5�R,*�W̡wvf������G�G}D�y�0PR���xf����h>�IO�8�	/0�C�����q\�ӳ�!
\z�/P1�yo�N�)2NUt����3ņ�{Ӑ�dGvE1�c�ɩ��
����}���M���7n�p��2^'s*����GZL�� u�F͎�V:�sdl��8�q��>�ۅ���~�獂�0zB�c���^�q���K'��U�b!d6�4}C^L�@�,qf��DQ��<�SI-	H�_�n Br ͺ�5�w"KH�n��E�S����[��;�ŨA����S#��eZ��d�
I�@^;���b��|��4�!;�P {����l$~"t���R��5 �d�uL
�nb��f>Y;�0�^q|���g:u��,S�0o�BG����B)b���p�@�����R��/DV��j=s����(��QL�ͼr�{{�pCᮠq�_�L��P��-��g�b �p1�y���»?���AwY��>�h����e{�,y�{�k>�gó"Z	����

�qd��<<Ș��z�ںY���W��W�}֊ꦉ������t�W�O���(zIc�~��O'��R0�1��
��X�j�_�Z�X���C��W�A�R��]�gF�<a����,bB� bs�%�3�phk���VM�oќ�-�vR���M��^d�c[�]ϰ,~P A�jq�sW�����P �ӧ S#ߊF��J��&qk*��䗨� \^���B�����#����f"^2�h�{`M�<�7�oaB&���|Q�d��1�K�E|W�.֟������?�������펕��XS
>���%�� �J!~2���P�$~�����2 �H���z��՛B�v;��xm�X�7k�C�n�h4�)2h,�}�*�ɭ1kHa���-'N�h�}x�x�}�`$��w���5~ĠS��!�`4�FXlxVHYEB    fa00    1e30MSo�}4�G[�~��3�\	�>�S��.*LU�q+%�G���Ur�^�>XM,Z},?����������CS_.�6s���)-=��Փ+�G&�wZ�ڶ~F�`�%J�K�>��Y4��NԠzՖ��u�V���VUϔ)o�Ҥ�w��o��;_ͩS>&�~��]��)�!��ʦ�3���g�E^�.mX�q�Ae�0�b��������k$s�M'w��R�ؼo��FV���Q<z��j,�� ax����� !O\D���b���X�Ri���,);t({%���z�����
O  D�-�o��^������_ox������`����@����KF�v-4ܩXgx�r��Ҿi� �d3]�#�M8��sXe��.1P�8�!v�u�5�i��;K��ie�-t����ޥѶ���� W�/��P.��y���� 0����s�C�	�L�����?�N2�����UB�Ԇ���{���mY�I�w%���	T�p�M��E�v=���k�&*����5�����2��ꍵ�q��b����f>(�dϥ�!V|N#�k���<��l��V�(B�c	{ X����]I�&�	��6� �D�LFb��LG��f�R�Ug`��Y:�gɞ���-S���
�n�R'�YJ�+Ǫ�x��dnf�@1	��S} U���x �C el�D�E�3��D�$��r�}h�^����j+�~��j��!ׁ-�����:�`�K�`��
K}�~��$t>7�	j��зM�J�]�p+רf�PE��Hv
skԟ���h
͕ J�������F�j^��7�L�*M�Q�Z�\��Z�O��������r��E�P��!M�fG|��'�Ŕ����L2�Ǽ�I�s=�W���]�֓/�!����c��I�����>�3J��0��fF{�`������3G|�>�z%!�ܕ�Dz �Oa>Ca)�SJ*�ZC�#�G�XJ�(��@-�7֯6
�P�+��,]qT�w	�,%*r�G6��K\ֹG4������lC.H�`����&��9�
:��-��!	���Z`�nCIE.��jB2L)�z��=�]J��#%��v{�
�FM�vHQËI~����z�rw��� �JϘnX���H�j�4)�ԕ��!��/��_�\[��S���U�5�:Ve}r��$\4�u��.�`w���I*"��)�����뿑�1��H�C��L5V+�v���^Y
ǹS�O������+���S��}�\i!���½��������*�>��Ok�������RLJ>���^LQ��cu�1�~�{�����XG�66��D��Zj�ˈ�A�%���%_-i ϯ��I�:�ذ�2twVd̈�tC��{�5��j���K�����k��S-�`�A�yVE�5��X����H>)��n>6��+3XDZ����B��!��5��/U�62�B�Fm�V��C�R��2XÛM��J x#���q���H�C��t/O	19������J�G�@�jSe�;����l��Jä��z{���g�#��R���Aw6fn����9��`ڤ�Q�#:2��m�(:jxн2Q�5��âVȅ_N|�*N& ɫ�d�ݾ�#�]:�5�C����:M m6X0���'�8܏ó�J���Xv��Ӓy�إ��v1)rr��K���TE@�I����0 ecM\4�����ɠ�GPe@�9A��ɔF�"{Z2����%�
 �iލD6�Y�k�xF�hds��3O��9� �e����ӫL�W�9�s���f��`�,UM���T�tm FZ��*̥b2������%�:[0���Ǭ�^L�8���s{�Fj.��dٷ�9>=If&�jT����d��Y
 Uk��&�(VP���"���_v_� ��K�6���k���c�GQ��O�WS��jr���n'kHGZC�%8l���ؽ�6��n��G�Q,h��Fwn��_N��i����dE�=�D��8췿�v�D|;#�7��9�@�������`D�}�Р� �K���)���dɅ2�[��Eur2��vv�*i�%��F �n�� �g�Z�jZij%����NO\��-�[�PN�J�.j��a��V��W�Y0�g����y蓶d���Z��$���6č"�-�f�1���~<��@Vݬ�u�\k�(�U"m΍w����^�i�b}�?�D��*:C�����H��m�9i}E=,a vw���Cvd�e�6&i����Ő5����h1�C�qc�QSm��<`�����OG���p�]d�~��l٣�������sD�P��C���g��� rǘ���a�o���Y��QtU�{�U���@�0X.�=��`��SOL,n���5��6�	��ֆu8D]�H������X�!��i� s��B�(emq��R��y^t):a#G�6�3	{�=#��\Z2��u�U���B�"C�L�g�xBzʒ�f�t�2q6�xE�V@p�F�FD1ο�3��('�V6(����l��M�ʠ��{��z�$���G�8�~������7
�~�v��W�bѧ��3���tH�R���b�m�6��^a�w�}Gc���(7��5�9��)�vn�*OP|���T-�MM`�8�J����`ck=��ӂB���_v\�Qƭ��zx������P\uF��B:�n��9��Dn�o�*1ECD�n���nc�k(���`���>2Z��`��p=4Da�'�-��3?ן����k.u��=��\�4R�/���z��M~�<��L7��i5GnPA*���L��W���`6�*Z�L�%���"h��1�Tv��R���z��X�־�mA��*��J�U��<�l�TP��s���U�w4R/�f= �ْ���=н�Qr�,#��S]2̱��Y����0|n�s�5�W�N��lx1�|c����L,w&"-��?��u�rȿR���m���卭��t�b�%w[�1�$����D�j
��8�ۿI��h[Dom ��l�-��	^�WbD����^��1h���I��/>]*��@�\��D.��fвp���wS���a��O�����v��l��������7�]	H�yI;ѝ�SD��L"-J��s;�>�='%��5B�@''�ܪƼ���/S���|1��FN/:���^ĀN��㊉�n�@]��]0�(KVko|~���e!&���h��%[���MZ�1�#��i$h�h���S�e�5+��|ޭ��rIJ�8��ob��c�0��9��?��q��ŻS��:�1*^��p3J��\Ëb� =`"��w�7�4c�Ő�v�m]����)?~g`��O?35b��N�*��P����|�C7����*�0N�މ��Ϫ�7!�]�<?K Yo��?;r��N�����,��Ӿ��ڛ|���&����Vخ���X�W��}μ0&S�-�8/ٌ&7���-���BV�Vz��쳢\��L�[q}�߬��A�y#{_��Ic�4c����8~�a�@�57���ς��)��Mi�����*���m�P�IW�%@�����F옆�#�-�?k�k�`�4��`,:׉��>{�2�A�s����#	�� �g�h�w�Ң~���Aѧ/��AAt�P�ו�Ů�Hm�����)ڀ���'����۪�r9[Rh�.�c0��̫�%�eʍ�
�9+���J��߻��A��}��՝q����jЂ�w�����&+��S�Ϣ<���Ԃ��8wg�1Š"���&+&Qlr�yZB�{ ��X��2��ۦ�0��J��χ�H�G���i	�7D/����'�U���Rɥa�E��[�{�u˻ۄ4���D=Q����	k�4�e�2|C6��52`#A���Z����n����c:dB��N�w9[p���aI�3rǂ���N���ŻlV��5~�Ӂ=D`T3f�A�[�גΈ%iąa!5S
�*��0͂�B��M{{��6zƇ��vXL$E&�����u��7�CK�����n0���zc@�d�����2� �(�깸1OR<a_/�`����xl<
��X��v�	������}H<Č�\[ne��#22�IM�bҁ��}� )��0�C+�$����X �]�
615K���0��S�,�R��B�H�z�?P8Pa2L���"^�)�����U^��Q<G����/����^JvXs�!b��=l鋵Q�֗sÐ���s��54b#<�O��;4�<G�������S X��p�_��w<y ��/�Z�I�ɩ��E��j��S��/�4�
{�G��;�f�XJ�����uު�LH�K�X���r囫�E=�Rn{�-�QvZ|��E�q��^�\�1�����k�\u��/]�X�g̽����!@J�
`��/�I��� r�%��Z�l�*���t��A@6�7���7����YZ�u�}�-��t^	����)���b����s-+O���t��֟���ʸ=hb^	��|'���>5�Nm�݃*r[�	M�=e&���'�1�ÀoHW#B�?�@�<[��y�~��L�n���PY��7���R�}Nk; eTc��U�T�穭qg��}4��`"	Qs�<ٽ,t�&���[Dݙ��o��U�]6"����7z����]��Y��~��w�=�����#�!K�7R8<ȧ�P��	�F̓��kʎ���k*��N>[H��̢2���>������/�Is�-���9�����'���糕��m�).|��]�6��C�@/8�k B"<Z?K$,�}���d�"�U �t�4C�2�4n3�\m4>�ƌ��eHǢ�6�����^�i�����)X�ԦI57�У
xB�ͱG���S6U��xU T@���࿒�Jֲo,��ޅ�!3�=����Y�pj��#�2'K���sß�c0š��I�e�n��l�|�et����!Y�w�}� [{M��Ŗ�t8}	+��h�j����A�{[����B@;W# ����_�1E��,e2�4&v�D�r��qg�Ղ��=z�\S�y�-v>g +zb��X,�NE4ec�t7�M����ZdS�}�	�-T�&6w"����~���&Y0ų�f_�������Lh�.Xf�	P<J/�D�>U�`iՕ~)4�7"�w|3�AM�,�f[r��C@�� ���4ܝ��������?�E�_�\D�*�.Y)���u�[�ڄ+����v,C�1�$&�4��~�!{O���=TK��M�g��͖B����h��(ZiO�Њ�k�`����;�Y�����-�;��l�b��}��<4���}�ъ��7�A��(�-FB������<�4�T���bT�Ǐ���rQʭG'_��Xf�ܳe<Sа�[�KֺH� �p��K�l��e�1��1�d�������#ϔb�q�i����?YUח�%T?�v�ǿ�"�79��Ĝ'��U۠��pe1W"��";����9�w�A�8�,�X��9*�}ԗG�%��m�_�^(����oD��|��rF.K��S+�}�W̆�V6.?�DU�N�)��T⮎D1餒�C��x8�&{��nS�A��Y���;'GLZ�W҇�	��fuO���M�h��_��m#��6A FP�^z���.��5��^��w�*A��V�7�����\�hZ��ʔ$'sb��I=�#��,Gx�hLZV���pf{.kޱ�\E��Q�������)+Fu-��J�&�2?�+^{�y���_���'&�ZY�C�%.��,tX�d)�%�-�#/(#�p���*�[=�F!�Čj�$�ĕ�f���}��ED�M����Y����3;�!�a<�QþZ�a��(M�ۢ�`��ʓ�H��"�G�A7���E�d˪F��&����_\�)ڔ|V�ޟ��:]iOD���a�	��-'c���6Ke�De�@F�)�)!����@UO�vɂ�����G�`:<�Ұ~ms��*�_M݊��o��P���r�0��|��}_��=��������ǥ
���k�~|A�l�-�»�����^���]?�Є21���v2ۄ�0,@+Iģ0�I��x��c�:�bS�<@���r5��m^\�&�������'������t��"�#�rKG+#�G�?!���58��i)jH�=3��%a?(�1qx�x]=�9�ɋ�̯��� \s-�E�:Y�~2/�r��i�J1+rU2��	#uP�c����Z9�?�d.4Ks��ԑk!6f�����f� �{5��-6A�U��8U�jU^��رC٢����U37vC.�@��w�$��B��?1�i��;�'S��*2��A��8��>1�W^��[�g����T�=�H<��}�_V��٩~Z�:J��J
d�SI�y����jz�I�W��s�q��nL7VBlDb�э`�-��Nx�Bt��);�a�lfd13���a|eH�0�vv�1���$*i!�i�	�����Nmo�-�T՗�d��a.Y�PUM��l~��E_
�ϕ�%�?P��|vEW����]GK9�n����f`%���V�Б���E(���a}1<C�������9����!��൸�_���;`�wZ� Ȓ�Ū`4�2�[ⶫ"��BfK�5�U�:���H������݇��4�JuTA�Ý�^%��[�#~D�ĿK�d�X>����4t)�j4.�J������Mm<��tkPhly�����X �P0:�֝^6�~N:��v1�,�E#gg&~���%4�F���������K�ks��YY��g6�t�|z�v�5�Ӂ�"���h��^���D�=Qow�����G��H�#r��1�Rg�6�m6j�?��2��e^p?	��q�4k��n�Ԏ2<�wǕ�=��,0���OV�hOC˩k~ ��OT�`$uM�ha.��ܟ�r��!n� �`z��p	 '��G��YY���?�����9�`�kF��6ζc��z�9�cڛ�Ϡ�Dp�=�s��	W�ll������]�Ej���(����d ��8�x�&��1�#j��Ûhu,�a�����ŻQ�@�
�!m��}4-�����1tB|fQ�Mh�Q���U+���Y(BC��w�Q� ��̑�R�_0�z���c9��e'��e.��³L)�奦d�_8(�(;nh�d���W�N���0�aH1��2��Cq�X�,�3�e�=�p��L�t<p�b�!C�hG+[|"2��۹����M��	�_7A�g�770y����U�m����=��Ӑ� ,�zg�+�E�Z?�ͼX';����A# �7�A�����@Ʋb��ۼZ<u�4�!=u�G��A�(��f���y�S��(Fv�mg�W�ܾ�e8K�.��k��><hu�ٌ�	��tv�Ǥ�n�0UC��	���ӫE�l�����fiʹɗ����`_�UDx߂ �/���N�~���f�Ni�2�k���o�mg^	~!�O:��+%l��M�sX(��[S�\�S�;!��y6�y�K�~��Oô��F�b���먽�{������QF'�M�1��E\�����E	 ?�C�/}�b9��
XlxVHYEB    fa00    1d20�OgZ�9�Kda�P��q���\e���iUe�}x�1|{Z��	�Iԏ{�/����v{�&[��v�5fz�"� ����2 �l�p��f
�c��Oɝ�TVe��5�PA�L�x���_=�5dT9���Ң��.#�bݏ���c[�y�5夶�|���&Ժ�SH�k#^V=] _�
|�9D \�){��
�#�������+̫��ӫ���w�<��2��*�C`5����N�$��\ᢶJ��,mi�����y��l�O��Q�B8K�rPΚBI��Uu����K
3���q�D��{IH7;�nT�%�}6��ݧ7�>�W��uz�/�W��doF�0��H���T�B"��KT���:'�`U@�K����Dގ	�0R��/�����i��2���8�p!6�H�Ʀ��s���>��� �����l9�>,O:�����#�C��ߞj��HBi�a/[�@�T^��J�,�>�"�s��{nW�EU��<#���k%������QY���}i������Q�*���70{Dɲv�93)*�3�)4�ig���n��Ze�%�$���V ����u��x{��9�R�@�6b+ű��2o6�x�ܱ�����ԯ ݻ>��f�v���5��3;�_#�?�2UZ;<�橀Ht��P`�!��j[,V	t ��Q�%��G�Ε;{���y�_ɡ�l�����O�{'���SmHx��;[1�U��Rh�
Mhp�^Y�� �:�5*�����í1�{�G�{C{̙J�I�a#��%,�Z����y����fx�f�eN�'�����5�Kk�|2��f�"A�m>��I��H'�w�<?� !l�Ƙw���L�
-;е;=�:�C6r�H�t�	lHRh/�&fo�~�yߺ��f��#e�8�r�2ӗ�����v��n5}S�מ[b���;��":��aҫ�_0�k��W%Μπ���=?U�*; �����B�7��ꉊ�b�mK��#���d�OQBo|��?�'�u�2����,��Ao�N�΢� 8�s��c����4���C��N`���<��J�Zv�y�%�L}VO��*ۤ)��L>��-�H1�:����mr�&�Z�Cx�~S�*���G�5M���Y�ø9/�(W��d_^�����.GQ}ͩ��CE�#��W�ꆀ�w)Y�j��T[�Pּ�������
:���@���sn�"�?%��:ks�r�o��p;�k֠$8�:�7@v�3�%�U���A����չ�ա,���gX�
���`�F�YѪ�۔�ݎbt��ܿ��������(�U0TF���ZN���#��k���GѦζ���J�o\O������f�o�#�\O����0�sX�dV�v ��<2�~51���2�(��7���˶@�2c��
j�7��	��\bj��B�-��A��=�k�(��m[��mv^j��>�L4�u��TWZ3��|�0���ݼ&���O�L��ֵ��-�����M�C��MΓ5�X3��f����&��V ~�&���� �-�t�C�����l:E}���"ߢ�.�Ns�;�`]��l��X�d:�&6�8ȴ�4�|]]5� �&�E��M��q�@�n��EA��I ˴���0�X���Ԟu����MD?���	�q�GWw��1��m�]ȧ$r��ē��+M$�)��:�+'rE�w����C_�<�<��5�-x�S�;=�f}oh�����$�{==0�b_�ncjc�B�M�g�R�[���Ҵ,��<=ZH����+6�0@0�<����RD6�Z�����K��}M�c&E�.c��Y�xaZ]��� �p�#���Z_,�=(hj����uZ4��|e�����١tB$\���I%�g2�E�Uc�t+��a�42�V���IW��B��%	uV������G^hw���"�d�!D�̱��w�!�Y[ndFH]A����=�1��M	��B[=^��Z�W��a|"��n��.amH�7/y�eu�HҺ�5 �sގ���I��G�fK���Vڔ��a�v7����E)�,��A�Z�>r�*��$*���$]�?"Aq�q�:�S^�3��Xwd4���ڝ4���a�[����pl^���1N_�О��a�,!��m��B�a�D�͗j|ռ-.���l�"}9����Χ
���?�qca�^{X6�0����}~ܦIo���.H�{i�@`���-bvig�r�K���l�J7S�b����%��5�#��d��̖����य़`�&<M�����{���Sa��v�q*km��^������E'�[�I�!�E����~
K`��s�9g}Pf׶����d66�,��R�5(1&�p�Jx�+ȟ��t�X���;�r LI�����C�x=s�����z|(v�B<�a�2ݱ�/�� ��{Ŋ`פ�+���q��ڙ�ͯ%��c�{�	L�e����3$P�-��E����ztm��*�\}l.$e�%s/���0��3/�h3"��^�k6�B*TP�N��@l��X�y��٥Q�e�A��k�B�y%ℒ�PN�[�F/8N6	�DiW�T���"n�dƘ�l�����g�W<�2ŕG��ה�Tg��f$���b 5z�g�؄mB�kY҄Lx<v�u0���SMXa�`U�8C�����3AX�+�W��l&�.�ϲ�:� �����&Ks?�I�?��)𹯭��iOj��}����N�/�ȝ��w ���3�E%2w�XJ�\�BNkTo��� �q��T�bde|+��nTsi��6�������*ԛ%阋I�1��U��^�]ڰ;��0��&Nn�be��D�
?ԝ#Ø(�e�����b`�������~�_�]4�csI�$2�1y.W�1&�q���C��`�=_�l;;�pNrf�K�α�M�e�qi0���)?��Y��}�J���U�/�ɧ�ے���3W���bk1�$- g��8�b�l�W�+�!-?��,"E�u�?.e�1�c}���߶�\�W��S޾b��H����־�x�gh��JA�ʼ��5Q��c�Z�:zcߡ��.����5�3 "�+��R-Eo�U��w�Q鸜Z�}�a�i��ХVa���h��N�P�h�0���8���Dk�����D��&ӥ�p>�>�
�8��%^]�+M�`�Er����Z`?D�q���*�3З2vUC�N]~|}
�r� �;\=����+T���ӿ��B �us���~Lc�A�j}Av�B�eM��q�|��|Srl6@�l���������lg~R����#�݃�nF�P��|��"b�X���d/�wT,�xU�ݎ�wB��x�>�Y��y�7�$��;2�M�r넣���x1��~����Op@1���n-C��2��l�;�$��Dh�>DI^��� �T�^���Ef>К���^~��TG� ��_���5�cQ�����[��V�򼖲q� �A%#ҳw����[�,&���c���ӈ�d��t���Q1��(���Z���7k�T��%���6�d�2�B{ۘQ]�vߙ[�k	��t���� X��Lxm�����u����iOu�l�}���^��1s>w�����-�*A�ȵ��w@�*�Y��^��Z80F��G���&9�SP�K�C��M��ˮ1�m���h{9p]}@�p���u��������q��:�%�A+>d6X�D
]VR��\�?�$������IO3�b�J�!�`���2����{#���);^1���f�1�f+��(d�/��K�]�K�(1XE�=բ9�ƣ�X��{��@ı�"-L�TÒ�><��$&�n�IVU�X^fW���m��}.�0E��G�V����t"�� WL�H2Kgoe�=k�ǀOްj��+qP�&ૹ�j����	3�|	�0�*2+�I��.\�z:����N�-�o�k��l,�'���ܮ,-�>�''�k�����R �&Y&���/�V����qR���f��$�1���tg�I��I΅�מOf��Ӳ*�i���*�*-������ Y��Q���<�I"��bt��Ed?���2m��<�&�������yf�8�n*����H�R��jK��Z�0D�w����(mH���_dM��sC^}�>��¡�Wɟ��� LQ�}_�Z�0���4����#����(P����� �VV���eq���� j�ϰ�Ë,��h��u%z���ߺZ��0�p&���=�=��#�$$,Fne�6��)�ʣ�{hQ������m��c���Jh�Rߺ>��e�H��9ɉZ{�^T�/v�f�P�Y���7x�i�aes�y��	��e#CUN߼�L ��b�|�uRnou\X�݆��m�̮���⢁6�'�da�2l�/�!\J��UQs
�U4]���F��}�`�x���3�����%�g������� Pu�����r�R��?��1������{#?��7�fUeH���Xe��F��R�x�z���!v�Ĝ��u�������ϔŃ+<n9m�[��L�bmb07�e]\p
`�,��a��=��X�"
�y�NY��|1yU��FWFN73�㜒���}�h���Y�5䭥�i�����)�Q{�U<�@���i��E]�Y�thO�J���*˕�����f}C׌M����czu����������E
O�i�8�.�Q��貅pŵ���H ��!�>&�!�U��M"|jHe�����c�]�S��7�ae}5��	֝�;���w$���btiȘ�r�->' ��Ǽ`����"�`�/ ��o�0��M�o�Q��oD2n� j%1F��v���2�_Op���F8҇H�ᐮI�[@t+��n��`�ۤ��JT�f��11{F�d�<��#�����6`�[7ĢL�㮫��������F7�X0���*����d��>;�U͑��f:LCF�a��P��tZFړ�ՠ41V��U���I���ߋ�
��'e	��=1j:l�,)p`��&U���]R[�=�p���0���T�W��#H;KK峛�y�|�B���H�D����C���[��=�}c�ȴ3�Jxþ����M�Z��aх5��=�Ϻ���qa�������A��ai�̊:��f���|��Z�n?ߤ�_K���Ap%*��#&l�����tv:6д�Z3+;=���0���(���K��WR{��Z�ڄտ��rޣwO�����֘�EC�������Ʈ���~���=�����~]�5L�`��*��I�{N��� ;�`��{іچw����KD��'�
����������WO7础���ˑb��{|��y0
���@���v�k�dTHoH��qH7�}��סk�2�%@�<�g�aS���/vwG>A �UYb��
0E��D�j����ԓ�KP�K��jH&A
�*.g�h��d��m�ZA�WV�$���)���󪔧Kk����X��6����gţ8<hϢъnU
~�X��0`���^%���0x�ܽ%��o��X�� m�}��T���`�/�P�Þ\!$���%g�Z*�č6��ukO�s��t��J�a��7���J)=<��-d��]d��D�-�q����5����VZN�k�G՛��� ��wW1�%��̝rz_^%6��[�v�zZϨAld�M��:��pX;�uэ�S�ǁ0v�б���G����[o�3�����-?�'�~u�C�+�/��+�a���G���
QO����u������~(��َ��k����-c�̢�I��vp�T�\��А�]%zbaѢE@�F�_�-a]��<5(v��ڕ�3���B����y9�P�E��=��H��M�۫x�a������p ��Z��/L�?t#�B,��w���h�_Jj��2�zӻ����3�;=±��	lt����R�-VD:�+�O��0:?`z}���%K�V-4o��v2��~Xı�K)˧S�5Y��.Gn&g��tl-D#vs5�9]�����`�ܩ�u����G/�GNGǑ�?!,�8\j�����v|'oS���k���?�k���1�NJZ��W�[:�Iޒv��41T��f�I����kB�On�,�J��Է�jm�?�1a�Y�?�d���W�+�9�|��4�~8 � ��v�lrdG�Y����4��D����p��$Ş��<�Bi��ٗ��c�a:� �U��HUgUH:
�u��/�ɲt�(�$ � �e��=~(9��������,s[O�\��0I�8X8�ȓO��P.ە\�* �6u&ABW��t����7��=З���H�/�c�WI�s�f��f妡��}��Gxd�B!BuU~�"��~�-dUjg���1b��u`�����2ꑤ��G�cx�7ۖ���;�V�:��TR[��=n�#���K���"�� ��pR���I���T�>���k~��S�W�%�=1|W���4L �%�T�|�D<���h�O���0b!A ¢|�/4G�#Z!�=(W�y�nP��wE��q<���m_��Nץ$�a;����}�'���P�9�n6Xz,�?�߄m��-��[��4�+
��',�;C>d�j�<�Z���q&��<�t�dQ�A��+��c� ��i��v��q�Q�?�Q�F�Y.����`$F���0Wy�o�O�eҥ�����N���Vz��:�,E:Q���N{v�$��a���S����t�Ö����u�4���X^�6	�j�V�*�8Δ�*���ϒA&�V^~!)�]3|��ai���_�s�n}D�h��{���T1�	�)N�	��^W�Ґt#ѕ���6V?s���2�9�$=����e97�N؜}�"�>s(�c��2ͩ�q��u��6�~�UU�U9 ���NYqCC~�\B�;q�y� )mkΆ�u���Y����x��"p�&JUܢr�|7~ۅM|�`��1�Pt��ܐ���2s��K�sׁ��M������	�ݍ�0���t�l�|nl��F2W1�Q Ӽg`�~�KO5�$��Qm q]�6�%�f����ڶ2��^b��#�͔� Dm�JX�M���qzf�ւ����X\G��.�Ĩ�Ja>�����D�N<x7�[�׽�2`O>�S`������� Ϣ�%�Kw��ڵ}���n����F��̵��AY�:�ݤ�S#G@"�6�1k�Pc��h�#ŵ�|Bճ�G��"���������<\z"a�v��,av������p�:�>oK�'�<��|���(u7�@�~��K�
�4�G�4ҬXlxVHYEB    fa00    1e20�٩�K��3���X�L�9g�j�!#=�~.�y~(p�@y~ݬ��
�<�#�٣�bo:�_�w~��?s�\�7:���'$��S~��i��^��\Y�����s�z����V���]��}]�+ D(�p Qz~�r���j��C0� D���q�`�\e��Z�,�q�`K�i�tk�=��O�|���SD��^��[��T}�ۯ�W�����t�l��@�S�%�����*36�c�i.U��r��/�Hÿ��SaP:�ڐ6����;�bi�<��M�Ѓ�Y�&�(����Lpԯ���Vv�;ĥ�FZJ�}���  ԩm1�婡X�#W��6�l?nו	���	���N��)U4���ئp�;�vY`�~֑L��Ki�a�a��XX<�4��A��*���	�f7��4�C!�;uG)Lf	�}�<�X���9��Bu����)���=8������؏1��i���bs�2ۍ�;ɛR��E�%�]�d���o���M��0��뫽�-�h�j�$�|�����>�z	y��QDo��h���4��+:�׸k��ݢ�5�K�-�)��P�ʜ�gLb���?�M+�է��̕�..n�A;o����[�c��m��~�ߓ(g�ܻk�~Ƕ09mNI�A��\� �Il/���,d� �C�Ȼ%[���ݤ���A���Ş����z�Zr�(���N�2�H�NӯA!��)^�����O3	"y'��K�R���ȠL���Qz:b��׮	ݓD��_���5Hv!��/P��d�C
ȲM���Nz�xւ�t���R4�2�VS�^��湏� ~_��୸eIF/=P-��~)�0�qh/v�H|zT"@�����󰚽�lϫ������4��9-�/s�����`���~�-s��� ��u�
&+��� ;�&�W�5X��&M�|q�7�m������I��I�Bq��C`����#Ոҭy�j�'�V�Z�S��Ex�< Vз�1�Vҙ��
![7�j�l��I�Z'����e�����4���;�9 �@kD����Ʃ�[$[��Y�����?���}��!�a�i�E��S��'d7���<U� ��d�A��h��F��HXl�/&�aL=iXkN��b�}%�uB�Ί��(�;�0������QJ�~|T��nON4wKD@��&e��
��9dd|����SL�ga��j(8��xq顫�!E;�GHv��O�YMN"�LGE(H`N�1�j�|)E�PeB�N��1��!��S=MɄuaa?"eM
��	�_��)��5���.��Lo3�*���1'�dpz��v����a̶D8�8�q"�ײ��K6'��+[�B�O��Ec���OfCVZ�F�v����Hy�i=������o7|�^w��Ԩ����05T_�F�m��]�T��{�Op��K���c��}.3��A�C��-�N�����b+r=#�W���_a�ś�蒛��j�r˟�rJ�YW��$%���R��K��z]Ҕ,�A��+�0��IbUeF3�K���P���zzsB8ݓ�,[�X?�L�C0��������8�ߢ���@���7�m��A@�Z�Xf�T\�d��/I�܅��е��U��q����;�a�yz��z�|P V#mwψ@��S$��@t�?%�ЧGe��cS��:�'�����w[����]f�����7ԣ[�����1a��ֿwC�!�78,g�D^S�,�'N5�R/i8lXG4��{	ˋ��q�P��d촵���@�� @��n�L��e�� �m���mr�{k������p6�ixA\��j/�ط�2�{�M��:��P��[� "�r
���cA�Ԛ�H%^�o��!���Y��i�V�
��b�/�`�����2d��J髠�Ke��˛��H?����l�ξ�d�����ֵ���o/\��-�Mʍ���jL���$|�F|�8�i,���U�� ���w8J��=�7�SZ��u���Q/2�yܝ���UX�f�	��2+N��\6Ɋ>������b�p�!3��/�K�Rjzk!���t�&@��L7K���x��ϋɯ:"��y�.��k���ѳgs+<�c��[5�ox`����Gi�V�Z�`�znU��܄m	��^��)�ԔQI���u'��G�������!2�z��󎘫�D$�D-���e4�I{�@����m�ߦju$ւ������p14�}*Q�� ���� ų� G���-�s ��!����c+���r��"�� ��ʆ|b͓\�C5��N�Q�e�`��sɮ�d]�/����H���:v��'��O�O2R��,k�<��ss��Ÿ	d��[�Wn��z���;��a@�jCI��-��!���h�jJ�� 
`�/+�=:�'U&zR]����72�NvC�����W��a���n���`�o 7L�e��L�2�G��^�j������i�ەl�4�.�Z�&W
���V�E��;�[��]E�.�pEf9QO-����d��3HjW�L�'��jF���7���q3{�Y���41�_�����\Es/�ܔ�T��������ʦ`����lBaaƑM�F|�|]�����ACE��,�f��b����]m��x�+�1s�x$���%FQ��J=Q�C�V�k�kz=����"l�a��Q���=��}�b{}��5�^�?��������������e�fA�����&������"��|Xj�@(�ݝ�3х��I�u�ۣ�o$Jl�&��^�s:_6$�SN(b��]���H<�����WhO=�ĮXʿ�|t�X��_�v=O�[�P:c��Sݔ�W�w
c �,e� /Y�M���V��7����m�x@ʿ�1��r^��]["�3��F�p��26��]���ᥙ2)�d�:/�z�80�y<r&fD��l��B����Ir�՘|��1 �N6"Ի��L���w�4a�5������ ~ �.�W��2�c���9����J�`��F�����~wM�b j8!�*�E����e�E��L�;Y�}���;P�[�ex�D��]kf���4�������[�m[���C)56=���<���gTo-�Y�|twI�f$q�����ͽ��bA��%%��f����e�D��W��qLP���'S�i=ցnmVN����K*r�>������B�y�_�<��r��t�˶ݙ�+�%� ��S�%:6�'C�}J1���I�X�?�1�����~��
�ɮàB&�@ˎ��)W����\f���/�/��x�����|�	��|�mH�K�a"���fy�6�=t!E���f���ڭ&S�OY{	�������?���9DѰ��hu��}�p��B��\�Iԛ�F�
[i���r�K`S�Uf^�q��`�uU@�HV�!�7h��>*��<�"�]q)�'��d�,漫�M��RK�] 	� '�U���됍i��</�e��Ƅ�4,3�s}p�u`B����Ռ/<Cr��
��6�C���c۴5�ؤV��ğ�,8�ӱ��4�w��~+k��,��Z�`�u������ׄ]�"�����7A*���b�A�8�}�FG[��Ġn�5���3N������G��q����؜+�M��sR��5��n��>L^~>&X��l�[�`�@q�����!1�e��6�F���	Ouk���4$3��ײY��L�ʯ_s/�����k��Q��闤[��3�ì�5z�l��TЪC�E�rPxԓ�ފ�j�e�niA�sI�^�$��y��o�b��Â�0���&��Ð���7.�����G�B��6�p	�\`�O��>`)���a�BH	�q�#��ߌNpH5�H��0��x(Pz+�{�s1Iy�R���v�J��Hͽ����vY� Oq��L��G��T��#%Y�3��@��l���߹f�Q�jTգ����\�*�>�u�u"���,����\,}�1�;�I@N�^�
��Ղ处��2@�^��W��t���o/�U֮#^��1�JjY]v��dv^ם|ݓ�o��F8g���v�K��I���1γ��������^	��r���_6��:³�ҏ8��zBO�N� 3��Du�fo�� �l��_9����&�/l�F��8C�0T~R��"o��p�>S���\�����pd�~�i�ʘ�:�ʅ�k������i�����~�^s��xm0u��:w���M���φ�J��c��Gwy��>��4l����p-L��U pδ���!��0�z	�w�]���{�uG�������]���^x�IP.e�',Nu���f���dzWo�_�TV�a_!M�ӭ�6|���;�cu�?��带~�yf#)p����.Ed^>����=���;�s��4LƠC=���&k��l`UG3�����A[�xܶi}�1�IrDvXp�ņ6�m�?ۖ�<>�P�p��Q�aU���t���L�IW����5�EӒ�惧a��s�C��V�+׽���b���2�ݩ0�"/6s�@�<�4t�V��P�]�;t��Y�FCM����h��� {�*��F˚h��nm���ݜ�ݢ��(�4?�\��ݭ6r��U�?)oӡ��~Y�+b*)y���}�%�ѳ>p�Yp*�q��Z	+��K��g�z
n���V
�sz�\ 9� �Э��A� TI�?e�~�(=<�Y��=>�#/��0 _�������X���+_}�:�1�4/�.�8���'�_�9��@B���w=�.܏�`���Ǩ� k��+L��)��^ZұZc�t�j8����Uz���l�#Q:����v���kejPLw�:����� JnG������7j�l�b��jt. H��2�a�Ώt��a�H|'k�g�B����G�ɬ���m�n��XLj�3d�}ó��g"���~���05ޙ��B5cC\ŉ��������c����Ŋ��1��W�G�-����Vu"�����n�j�V�H ��;���>��U�mf%��������*\�T������`b��f��{쀷9	;f���������:Y��=ռ��R�<�����G'fе������x�s���v+�	pC���(XZ�7Ϭbs���5$�Ghq�0������ ���
C��[8�T�_�i���N(���@�L5��v���yX����9���Ar���Pe;�_=;Q�{n�������>$���}�[#�*�+��?�;�8HtE���?���JOp����T���N�/ڄ���X����P���*���ahnA�[ry�"Ʌo�~��tT�s*�т�]��T��J����5R�iռT����@�æo��Z�������u�6�����V�a�2��s�âf'^QV�����>c���F5�INZDxT2C]~K�:��6W��]0�I���8���6�߭o����:��G��,����?��ɷ�o��	G�{��ߌ(2���!��=�����ci
�� P�,�ܵ)���"����n�7����#$%{�e�m���R��	�
21�R
�b�ϰ/�������vĊ�]��_}h,z���[�{��[�#�k�b1o�����b̾HD�+�O���*�a���e���kV���>ky�f��_�O����Λ��<E������	��E%5)m�#y ��v�ٕܢ�j0�p��	]�g8�c�9c�
B�N����v���*��%�����G���Sl��_��w�����j  n�՜q�r�U���B�lw�;" �=�l��Q²���Q��h�Z��iLk�¤"�TDsr!��+=��,�b,�T���� ��o�����8	�Vk��+���OѮL�G͂�#���%�����QH��z~�}�{��m�sW����l�cV7و�8l���U�6�{��"v�o��)�[J!'?%?�4���)���:�NygxꨥG�M�F��S��K�0��� ��!�a���^��}����,�QfS���$;��^c4Wn1����8t�� -<#�*j��>��%B=���:ToPC�,i�|���~�.O�0i�{��R��m�C�K;�k�@����O�FSå���%�:���ǯ4^�;�#�T �Co|��|a� �����=���d|����d�#�J����ĵ\U�b��OjH2���ʠ��^@4{g}�I�����^m��u�"�1%�]N��5.�����/���M�-��Xk��%�_~(�	�F��[j���
�v˝���"���<��~�r7ṿX+�F4A�� w�7��ٌyvbyUD�ks��7a��x��A
�8ۃ�����*}�*?�χ�zT2-��ք�~��+���Y��e)��za� �Ǹ[�4�x�P��ѥ�0M��@Z0)��� �J@�/o��Q1�=��c���i
n����R�h���$���	��{�R��p�@ό���u)��@(e'zՏ��]�>I��l�{�*|[W������y�B{�|�.�v� 1l
�?���_�"n6Ҟ"�H'�a�u�Ÿ[k���0̒X��\'��2S;��pm\��"�~6�~����g�mg�����}{��0�u�l���PO�)8��-p#!�.\�4��t����[K����[n���Uѷet�{4��hSj�P�Õ�f���M����4s~�IK��}� ��;��2Ԓ���t^PM�՘���6���鞍a�[���傛[s�7�e�^���uv��&9�g?&���� `�Er>�m�.�_���M��@���m��)ِ��Mo�K��+�	��]�b`�*��P��A���������ȭ��m��P����H�E8y~�ߓhh�..{ǥ��S�0ϟ��pQ�8����$m��ds��v>�c��o#I���a�B������ц�O��'�_O��7E�D�m�ђA�~G*�|
�4��jdF!`�vP���e����]������-U�~a�Bz��zz5�0�����`H7Kщ�'��AފcCk=��ԏ�!�EH�1)z�OE&W�-*̢��}.���^���=������Fn�0����@���Y�Ov�P5��x�s�t��?��y9�$gy*��t�đ�V��������]�%|/<���UL�	�O�|#s��?|_�}O�uHP�<j�)�۱U�T���/���+������D�^��ZC�������P�<ƞ�q�|�t���>fJ���oi��[�i����7�˩�|�9�6�o��>�f_0{�K���&��Wl`%�m�έ�u {�T�j�B�|�L��,���g|��}�1�oRV�pK?n���I�@�3�'kth���o�_�N��,mh��VE��%ƍtķ#H�=�r�}.�8���z�`"0r�vUj���h�
�e����%�+��!��O�b�H���N��_�Rl�1� ����1Pw~��]`�pY�\-d��g�@��&��ӈՍ����o�CG���.�>�d}ݲ�~�1Q��R7;���̅v�
ċcT��}Z�/��g��6����}i���U;�ܠ��'{h9��>E�g�����_�!xz�['���h��B�����wXlxVHYEB    fa00    1e50�%a���S���"KcDc��,��#/��u�4�q]4(���G��ɞ׏�0�{����~�8ؒ�9C���S�LްvR���UX?Y������YRf�FH�Z㮮���&9b�����J�H��-��TF�;D���=�Iߓ@4r3m��~O��xoFPVwj�vl��0^`l��B&z���5���u��Bj+�ʻ�]p�"q�\�!�Lc���a� ^�����c���0�,k��0*׊���?��NL�σ;Y��{�~�v-������M7s2��;�B�%(�p{O�r��M��J��NI�xs~_*�9��ʴZ��Y�4��f9	������N�kWO���XT�n=��;���4{��A�e�F��{��|HQm����(�r��{~�<��5�a�"�>uE$��r��$ mXDm��w���J�UU�3{��W��x%A��0.�/���@�X!г��������(N\��3���K:.�>:�`x�$�n1W����Dtb��
�����^C3��Z�
���Q�8!��4�(�6���󆹎��f`R)a3�6�Q»��Ě!�낾�+&�O��e�.<[V�m�,�3�0�HW�3��Wl�Tr��a����}-##�̱0��Ǚi~�J(4�iM3n���)0��M�ᰍK¬}&�sN� �lF����{lc�AS�|̀�?�jF�ǘCM[�"�]��x"O՘��9��Г� Qp�	�0�,M�G��j}���CWoU��(�tb#b ��3���e\�˰�i�d1RqdI}��r��@$e��?������BE(�!׷JG_N%��Qnڗ.�0��7�e��1i�K�D5��Lbmp�[��q��D��ŷ� ��T�@ b��\���S�:>8<5&�q��yr��T ��G׍�Kkf�FT��AD���
�2��з��C�v��wR��-��2�Hpd֯I����Y��[�妮Dek��aFdA�ێ�)G��1z�����؈�9�4����������y]S[E�)���0�y��W���/^�����V%���_@#m_��]0A�uO�5:^�W�;kF�B�/�b���7��D�WM�2�3`��c5���3s��w�+�-����&�5���1X
XW��Ӟ$��\��,'���t���֏=�?��1�U��_�
Զ�G�?�����O%dl�UP�����vܣa�}z&{��OhR������kC�����I=������Ӗ��m��C��+�F!�ߎ|��+����f��ۊ���ً����mv���~� � A��܈lp#��坽ȇf5_�n�8+���]֌�q����S���T�qnދ��CC�E�f�r���6~��,��c���HS�$S$6����+���!�t��gF�)pG=[/�a�V���.8�_���C?��}�@�t9�ë����#��k��/m��@�Ė5��GS�[b�,�������*�΅N4�R��?0����Q��K�������X�=UR:B����f�@��&N+�`��O
t��ގ~6�@���"�Eh�R{;RI<��N���'��z+��~o���7b�m��|�@�[��ɧcB}�Zp����(+�$z����G��-��%�Og��I�� \H�p|�P�Y�CJX����^�*���J�V��U��L��n��jp��UC�|j�J��������#���_��k��2�j3�mȨ�BQ-n�Zŧ��[��?�S����7��;g82C:!�(�@�$7I��g��n)t�����t*���I�g^t]�ZB2���j^��flF
3?ۖ��5�W�����'4���+	Co���6�u�}q��h-l�Jˑ(�\8U��r�'���r�$���������x|�'H�6�I�}��@��Z�o��mx!23�ޜu7z����7,����Mxk�m9O)�d�s*�T��>�Oa��Eu���bԖ�7�p�����
� �f�Y61�%�l@�!�2�+�;��@�!��$ �
7=��ې ?��RP��C` �}]�y	ky�<g�8��J^��p�u+�{��<�cކ&v���2 W�ѧ�2B'~
��D�9��Ź/�?
�bs|�_ܹ	!3<��9v�n��+�5�]$�۫#�x��(��jף6!�tESU��w;���ް	�s����wc��%� �3=A�6ia�� [t�Ĭ�`ɔ���DWTUƁ$�P���6W'Cr���Լ��	tkp�6������P�E!R�ѽt x,0L	�Ƈ@��a<����<6����@Q��c��)���͢\,�]�O���N�!K������u��<����k��cjPI�=��V����K���mSHu��?�%O�ȢN@�P|�l�n�#K�?����l���hN�0��I;j���P�%�C�#P�{� ����Ld�5!����0��QY8M`�\/��M�P�"W�1n��C;h�o%{>Р���?U;AŐ�=�M�Z��N%�?�t����RH��z���Qs0(?���CbL���p����0�ª����l
�	~�^���/%y�B��ȄF��� �M}	ȾƖ�����a���/զBe۷*���Z�u��h:WaC����:F� �}M$;i��z�b�����B����~{<m��	���'NH�Tw��n.�T�&�>����.}
���[����-ⱚL�I����k�jK�^�f�zit��w��y놹�& #���f��.O+����k�G�7u�N�K�2�,߶f�;Z���������LR}[�''����~~��R?R�7���_<ĸ+-� ��D"���]MӞ��<�mZ�Z;��o�����S�5�Ւ�X'�L�
\ߵz�ao"�	_1e^Jds��/�~VT��NwQ���P���a�K󦿿�w�'��؆�����+w0q��jw)���&��YX�0K%	��}_"u�"�����KQ�`��DT�J"�nܼ/�����_E�F�	"�A���R)�%��NU���H��p�-0�J*&�%�ѻ��}���ĢH��R1݋L�zx���6x�;w?��L��o�$$���|�iȸ0����~*�>����{	e^`Q�J��Ҽ�V�ܴ�kn](�������}���l�l�_8���KA��V����n7���5��+�0�ŏ��x����.J��A����^��h9����0�_�8U�����7��Z�Oę&�)�&��, ��@�yr+�gXX���*eU���ݐ�k'�(��*>���r�w]�u�w��Z/�<W)�Q}K��
�)!���K��ӧj5���0l�����gu�4Z�"����rC\N��zqk<<c�����ʙ��-�potDG��g�W��nA�x��~3��ҥ��p��,�6�%"O.7��������c!r��(5��!��C6o���VĜOAC���S,�>�d��g��TB�!�!�Mj��s":I��>F��y��ʳ\N@�UR6��>�:'�G-B�gQ���{9�m��	V�0	���o~���Ꟶ�12S��*�/��-�^J��K�
3�4@�#z�g�_�;��`A��=�tͯ6�Y��w��
%�u��oҟ����7�Љ/7v�~XQnAR�u?hU�����qH~���ndi5d,}d8N��a�o��T�խ{
�=��@I�I���v��|��FshvGM� }ꮏ���DlL1N�dl""��r��$R��d��P�'����5Lx��]��t���oՑ=K�q�
N #I���&���MF�
田&5�M�̘��Ոa݂ûF�9ު%�����1�s��R��̏���z]a�� LQ���y���,���B��l�P���ã��&��QO���L�����w�R�_��A�R#��δ�/r4w����Է�͍�.�' 8i@��&
�%�i؂��un��[���C�6E�j��o��K��̓�>B;.#��D�P[�ڞm���&ST��耰L*m/����/ʹ�ӯ��)�x�P}G{��H5�g����=�A�����|��pD��Ecm1�$Y������gL��fA�?���Kp������3?�����(��f�ڜ=���f��.�Y���\�O��0�4�O�@!y�����'�Nha�-^đ�-sKl���|�SM�/_K*�i�g'��g�e�����=�8���6�	�i�I��l�֛:k2���½(9lL��t	�����^�����Œ�W҆a���/u���P���tϙx�`B�w���|%d%@�ئc��b�Wb�U�e`1�~�z�o��WB���%b|U�%�O���Oj�Q�7�WE�S�ٰ�׻oG6&Md�L-a%����Wk��V���P?-����5E�m�թ�A+�A��z-򻓴⮏�G9F��G�lZl�j��j���KO��n��˷/� �q[�����r�4#�2���L��-L�2|��g5ΒW#�r� z�-=cIώD�\އN�h���� �.;��v��I�� e�}�,� �0ʐ��l��� �3↏����\\g���b���#( �φB��Ъ6���v)���k�Z��}d
��j�qi�����Վ�i1> �u�JѤ�ͦL�����.i�_�?BdH���L�û�� �,�&���E��2P�DHN�44�|���r���U�։8�"J�rc�*K��?｟�˴B�Ol8�nw�ޭ\� �ǫ���V��*��g��C,$�$zyt�� �W��a,H�VI,�|)��Wʑ�����H�9�?}���ėJk"��<���� �f{�x6�l�[fP��_������ߔ,�1�����U��l�W>�ocW��b���(�W�!�#�����@���m$����f:���9�@Kb䷰�/��aq�~�F[�dKfM������Ե�*����Sz������$qo���8�0�7�7+���y=F�y#;P����z�a��3/F�>L`"j����I�ZQ���ȉG(�%�u#�X�p��bkj6�c�:��'Ԩ�=�NB��2��*ή�U��J; �[�J�K]�\�%3�����$�5v���I?��q�(���l+^���$��NA�֥�!��)d��f���o"��c�y�|¿��s�]�f�Ug8O��>!q=Ħ&� G���}��M)�*� ��A��QlA�M粴Cw-�>6����R�J���1L���n�v��(��޺.%�I�}7���>��s�i�s�N�cʁ��1�M`Hnf� ��tG\��*�쀋au�3to�6����j{_4�����]�U�	�%�	yd����Q��zw��v��]��a���W):�}�,r{�p���^��E�	���S�mG�r`�{��K�h�ۭ|x��Ϳ��\QV��Vn�w!�7�K߷�$�U($b�_�_ߥ��
IP�`f�w� �V
k�uX�b����{�lCi��b[�=���}`� <���k8̭���FL���	��K���n�H�IQ���K(��ÏtRPS�-��^�5`)l�a�s��@}��zFl��() ��n���&��d��z�؊���S��T�~xN�H��n{I_�w���T��S sﱠ����og�įy�͑�:wD��E�Ĺi�ͽVu�$�n�+�0����5��o���Ĳ\j�^���,�D�x���:y�?I��G��6B���f��k���~8�WuK�>h�H߹�Z�^��Uz�}�r�7#[M�[�2�cw���~��R��'
��%)����aEIhZ|�H��7U��w��(�0�-�
���A�S��rJ�٥�p�1~�n���NpYN�iJ��n���@p�W���(�����X!��be;}��D6\���Q~Qm�I1���"Q�@�>�<���N��c9� ����B���w�8�"�1�@� �c��'��O�����>����j��L±'��1���i�	D�'�GݒI=Qkw�E�����zs��x�!Y����GO�º�3��4Ⱥ=����ΚIG��R�F� �$$�R�G�)����'�hԒѸ��N���;~Md����b	b�$����U)%�2��`%(A���	Η��9_*p6&F�p`�ݑn|?UZK��`��h���L�{�R(�`�*�����Ŏ�뗟k��hF�4z���r, !�V�N��㤍Zs`?��Fe�*$��uq��YֺL�/���e�z�B��gi�@"��d{���b������ȃ5�P<:�l�xzE����i�ϒ���k�e>��������"��v��o�M�a
Qu�� ��{��<�f���DaC���&<L؞�B�ZB��b�'���z�A���xA]hh�3�JY����6�G��ma9��-
�H�z>�e�]�����KBj#XvW}�P�:�&]]�m�XWr�i�}�6��\�U7%��ͨ��0�J���n<WEʛ�򧭪�]�c�J��[��� �I�w]��G㓇�tsy�n�
n�e��.թd���<P<�2�><ͫ���B|���#�I$=vl�-)��.���A�{b��H�� �'�9�Ml��"���m69@s��ʻ�Dό�[W+m�_�x�\daD����{6l�;�/��N@lG���h}�b������H���惬�ﶞk��C~@PB�����9�����q�q�Ij�/�!�艩�Ww��|����Ǻ�{�����|7(;3o��l�v�iYg<���vS����~=���ŀcQ(௢��s3������C�� aQ���I�j�dқ޶�K����P.��`,��;�x��|��<��wɡ������	rI�덬��m5~�G㹼���ZE�g�/K[���qt�a����{������=��pGf��e\��̲ c|���;;����vV_7\:-�0s��;36C������`Q�h���h�?���,�g>ތV������Y�k��RW���oղy.����BU� �B�����U,���=м⣞K�I��]���;X��\z�� ���&{����E���}l�ҵ���+��*�Ԍ��Y��%;�4��ڠp����ە��6��寖zr�$c�O�D��h0�,��:��ɌT��M7��m��NH�b�6%ˮ���.�h�+(�i�)�����s�S-�����)IF<�ɏz�Ö�L�9h�h���j�2!G�c��&�W �I7bT0�#r�R��0F7�����@�s|%�Y�����@�ET Z�^��.�'���$�ix��O�g�<����o �:�[���{��`j��LҨK����M��7��+��.�@�ư �~E%.;-R���@��	U�݇H5�5
c����hTݒ�8�q�Z����څ���j¨!G�q�~A����U3�F`��\'��|C���Nm!�� K�n�b��ө�u�.�+c ���*�C��I�淜���*�ٖt�,�*�����+�����,/B�?<5l�`l�S(0&	�#L_��R�T�.h#j�0X��:�8XlxVHYEB    fa00    1da0}��+�ʝ�Hp��5���{��҅VA�:E\k9���72C��E�Z�O�G�R��V�̼N�F%r�񎷣�2�=al�*�̗�����/TOe�����r�$>;�T* OP���K�;$"��D�0l��jw���'���i�W^T�tGN�Ta@�H����ِf����d8�,Ө�L�b(�zph�k�RǓ{�1ţƇG�g�\�vp��s���G��CH�ק���c'��<��[T{�ݵ����t8α�GbS���S{�B��1,��/�'a�	�u�A�Q�!$A�j˽��nx�5�N��E�����I��r����k,���s�g%�v��J*s=˟c:A����[�Y���h�b�9��u�ϻ Y�Ek�p�Z�-7�I����0+�i��q��W��8U�S��P�~3�+ר��c�o�F\��ض�r���gq%����h���-�ܯz��_��g��V�+��Ȏ�O�����.�����8�T?�p���Z��7;=�:b����o��OhI{��V�,��&��䟌�I�3u�����
��A��h\?��+�wD����9a��Ƃ1�(Q)���2)E����	& ��X��c�+m:^�a�vE"�S �жKM��H�����g�:"|��1B?���m=V��@n���O��5����h?�^A@������R>�I×�r��������omv���$?vP��A-i�g�x�vA�^m���)�	�F�����O8�m�K��	�ZQD XB4΃L�0=����1�^�
���'��*�T��o�o�|J0�E��M3�xn+�υ9(��8`7~
^���M���ܠ����E>S)�8�Tƫ�Л0��c���>>-)�W���� i�#�u��a(�mό'��>�6V�@��F��pd�~���̥Po1]g�]�P0����Q0����ϲ��l .4c!���9v�H�r:mD^�-���4���&ث�A��<��������O��A"���-�{�V7* i0��7�A����D�|?o�V�C�@fޫ�[,�Cݻqsc�Δ�����L�Gף��t�﷏�Ʈ�zʟ�C\E���H��ό}�Z1�^���?����KV!`�m�X���u4��Äg�߈�݊1���������N&�h�-J�8a$�Z+j��8���(�'�^~�_�i�Y@�^4u�7���� �(Q���5�th�#��m��`�]k�[l��)*HX��D��(I�r5�մIк��,��7�tO��Ev�j=�h�o�B�զ5#���Γ
�#H�/g5f����S���u�{�aw�gG��#�Q���,pN8iV5�c����ӷ��8��9"�
x�x�>�sQ^��^����{�?��=V�N.����z5�	> ?
�H1#�j��7��'@�1�%�/+� ��58��̾�;��&��� vm��q�@c��:����P��e�v'ipI���Rf2����*u�8��,#�2ǥ=���䬉Ee��S{�8`�Ĕ/�>�I����z���J{B�f44�;�����R��9nҩ ̜��拪r�U�s�╇�ld��dT�;FhS7K�z���ȇ0�۱�-�������9����A�����-"`�ql�~ŴL��a8�#�㓷u��9���^m�{I�G����E�~��}�k��7?�
������-��1lI']�ES9�k������>�O�Q�A����
���8B�鮞��I���;�bL��f���FնcI5!�w�Y���z�2��Sa<�]��"�zs�G���C
��X��|źpR})'�@�=kD��?ӂ*%��z+Wo�)F�+0f�9�Fhl�� ��32�?O 9��d�J�"�_i�Сmp�LI׼���|_�>�|���e �*Eo�����=HT)���;���f�(�a�T�-ս�)���El�я�8v}t��9 Q!�L���n���h�^$o˜�.����t)L���YyU������ڃX~Z�ǎ�ZOH��M�W�P¶4��3�����d�}|�	�d�0z�jk�{��c�KCU�q�� ���>lf�U[yKRj��L\��3��^���A���'�
�����Q��9,Bׯ�Ʀ������U4L��IN�x���B����g��E�Q�V\Q�3﫯����j�z�n��EK�qk�v#���VW��)�X�A���_A�+[�u�J��/Zy���/U�M���|V�|�m�
@V*M=��
���`Y*����x�J=��%��ج`��%[,�A����M���ޒoJ��b6����{ș���t��xކ�e��kOJ&X��"�_m�j[Fa
_�:�I�@-r
}V��
�݈0WP<�	Y�x����!�y�x�8 $n�?���2=��J�9�	^�5b�-v���Ȫ�=��.r���Bq>䒎�U�˶B�p��Y�Z-���q3b6p��A�mo��e��"�7��~����('��~��(d\o����W����mB�)-��/��2:dI��O�L�5b�3���C �1y����ysS��R_d@�C��Y�z�!�?_�A/���ێ^�!��V��҉�3�p��ƒP�^]��Gf�X��g���F[���O�ԉ�@{�		4P
��%])a�F�U�0A���}��#�f���l�鮞fm{��kM\�]HGy��U���cޥ��u����4�p�NA�gg����d���wR������:�K^��0��\Z�S���Ģ��$�c��$�X��O�udt3W���?H`�u��'�HU���>	�2فA���\��~�'ğXl��k���G�����w��,�����|q�5įv���Ĳ]z�X��1b����\�yN�߿�Y��v�i]�{·^3GEKF�@=k��wljA�Q�WX�C�!D�0;�� ��n}Րf�E+�7C8�^�M�xAښ ���t>�=
��q��y�ܹ���]9������џ�krc����W��"N�V�X�n�� x)��ӜL���W��qʫ�+���x6�i����V�^˒�ل�nQ�2t!��{������������g}`Rn��D�W,�^��>��	+�O���jeon��;	��ˊk�[)�«�%#�.���-^��E24�v	H�4�|Fe�y��M��zXF����Tc�qs�����-/�nΫ+��������\',�#0��Oa��K��FD-�9���<a�P��P�k�c{�`���g]�]�	Pk��*%��t�.�����F�	1��5��$�'"G �t��O��W�q�E3���4��f�E� ����E��^�(������SyY����%qb$�mv�O~_<�ܤ��!���8%Ӄ�3��oD���VԀ�i,@�\K4�������8�����C5<Gu�;Yy;�8^nr��Fr}�4q-tF�D�=Ts��d���m2�Фb7y��B���z�������w0�_���#5o�e)�k��~�b܇����S�� BH���;�����X<�J��Ϛ�[���ъK���^+^��8����ش��ݹR�Uo������ê��)��n۵\�ˤ=���O�� q����=Va[n���w�w#�q�J:"����� ;���S\��0��x)Rʽ`�.�{��OH)��j6�o�'���f+���*R��ix��2��ZqZ(��w�Y7߽�i�;�$!����=�.���7 �q�|��{yx����z�ZƑ`���K5k*lmf,ł<�+Sd�~��P�|���K�cZ:/b��j́�d�r�'��#3G�uim\�ǩ-+�͆y��(�+�V���(�"�
|�h���V6�T-��0	�h%a�\��`��#��=CZ4��L_B�|�ߓ9�J�Q%(�Mw��)C��|�z��j7��8�
e��H���XEO�P1鿸I\�!.��n��4B�����Q-��?�����o�����ӄ<VS����E?���)��ott��r)%�w�|<~�FGYwNQ���<��H�CcsG�b�3�:C�]
�ȸ�J��]^�ZJg^�'��d{t,J	�*�!�L����
����8Z5�Mt�%��M����cR	H����m�E>z�, p�2�ZRG���>AwRM�SmǭP�Wp�DH�Ѕ��w��٧r 5?@V�`V�!o�Yo�_���_%��o��S���,J����L�&5����/�:��p�h/F������QOL[�{�j���lސ����N�
x^�&<�l����Ń`J͇��l]t��Z�x
�b��������jB�z���T������R{��Y��zl^]�c9yo3s���,�(��d�$��c��'xEО)�������$<5CxR��S�aL�������=S�i�u���m^�Bϲ}�����]��-��W��;�D�߅*g���u���Ԙ�q��;���|�T48^޸��I��%�y��?�Y���p���J}R��2�3�(�j�uwy`��(O�Ӭ-��E�����O�M9��)J�{Fp>�ڟ��c��a�36����bmD�i�! X�Z�[�bfn����%� �f0OM�����P�4�wX:v�`c?`���L����:g^\2$�A(CH�綑�25��i?W��Hw,���R��RP��Ut�����w�Z���������@
�;BG�}*�����b�} }=.6��ØUi��X]%k���T��?�n�=�P����Ȉ�Þf����*��G��D��r(�0�E�A�竀,��]�������kƴv1���q��W��%�'���L��+\�nc�š=��GM�Y�j�0[��y�>�GL��<m� 	����WOiU����^@-R�M��.4�/Y��O�2j�{�#�<B^���õ1d�)4���?�
 �߼v�]N�\����v0�EZ�\�I� k�*R����b������z��P3����Y�ڨ���&_5 Κ2!9=[�3(-�������J����{[��oJڭ���Q˼��uV;�����6w����\9��Q���N)�u}�bU8��:~|:ʴ'ŁR����b�I� ��r�S���u$י|��&0��Xi����@���X`$J^	�|ق�ݗ�a����_*bm����׉��Dڕ��`�kXO&����@z�HŐ�@3$,�*�Gg�I h��N��Ə�@�2��vm%�Ft&Hmi����ȷɧ���O&�N;����-��[F�2	��|f�����]�3&S��j�,G���De�:V��<���g����3���S �|q��i=R��[�t���7����Ү~��.<$���%i���*��'Q�᫩�jD�:���s���+��.���k�eҟ�e�)c��Z��x�?�4����?E}^�'PQ4 ��
XmO�3��j��Dt�"�1��*n��D�İ��
��-���p��^�M�8����{F���K��㧛Rc��H��e���_;�k!�E�m�d��5Zu8Ý���� �P*����Q�������RȻ$V�, ߦ������K��*�ne��<���I��h��c��u���8�TE_�@U�������'�j��*^a�u���*c�o17F�� ��ݣ^�F�pLc�o5]\���݌� ����݆;wJmҷ�Z� m����uW��n�\uy���`�v)S�;�+�|��Z\���;�3JB�"T�1�RE39B[Ͼ���qh�E�77�˽�uuϸ��	C
y� �9�� �C��,�����c6�Ѥ�]�S��M!o��b�f�������ٱ�nRm\1�W���?�=��]��.<�P�+�u� ]h�,���X�.zބ�\i�ov1�|6i%͎���
��V��g��r��_��.]��)��q�����DM��h��	V{���#[�9����zͬ]�:\=�l���I�ΩZC/��0�K���F�WTB�y ���Ò#5���]r;Ҽ!>D҅�ch�7���l #�H��z��J9�j#��a�NP�Kooc�]�t3��-���N>����5$*�Ҟ{����,�G[���Ε e�����a�.3s���Yv��K]-���Sʸ'k���j���J_PL��t����|�uo[Hɻ�ng�R:�<��2����Ѐp��8]E� =dX/��Fm����\����/�0|
�N�f
���EJ��'|P��9�EΛ��Qབྷ��\����*�uU�����j%�����KPxby\�����0�N[JR**{��ǡ���aT�yM�'���i}>(�Ol��I�����H�$?����i*8����đ<V�aG��A�t.@Qc�I�L��-	][��C��\�����Hh%P�i�
�>LM�]ٲY�{�n[۷���\�?T�o�{��a��6��1Zs�(r��WƄ�e�� +�]g��˫V��1����D��;�o�8V,1f	�B��^΃j2��*)�cRY���W�W�eUt��`X�]Q�P�����y��#%n-ɝ��@�F���"N3.��9j�7���
Ǎ\�@(�do�:�J�B��N9񈋾K�F��Φ�
p����d���{��(+k�|�(����}+��V���a��0�ʻq-�]��@�v�����2/oz���E�p W�&���A��0WU�����A�~#Pjy;U&��l��h��l!�Vp7�j�GC��؁]�/���@������5!_���H����,��d ��J��$ Å+
ܡf�<pU�Xs"���ڼ�}�3oh��N�Yۍֶ�u`����s���1�'�#��^L�F$�,2:�u���8p�:<s7t����oU9y���S�C��x*���Q��_��d��+#Y&���r�B�'\す�|@,�3
�+������<ڳw�2�BN��t���]�����⟖�+��`g�ޗ��k����Q����fh>,@�y�6��_��ݚ��9��́�qP�R���,Pf���t���W�n��Q�[8�����!�n��������ӿDl�JM��q��Զ�,UxriJKMh�V��I�z�J��]tݾ�S3���F� F������8� !R_���xۈ#-�����Q�y9�!��F�I�>h+��~Hx�_`u���c���֝���|vgKNuV�91�!kǟ��pL�h��Y����a3�$��2Ǫ�r'�{h`����M!f����.^'���\�^q����� ��_������zq�H�f��V}ʠ�-�'[5Th�����Âm��5d��s�HO��G8\��������Z��'��uª+����-.g�+�����&[�]�h�9�$Ug\`�R���$aY��E�\�vOr����0�,��G�6,�XlxVHYEB    f314    1b50��A�`�N��
�Bۆ�휰w����̭a�3Ru�ٹ���d�̗�K�y?�ׄ�f�ԛJ�u$Z�|�����68S�E0M�5q9��~�:q�!'���%c��I�)i��@��J�̷ey�F��Wx���
�_'�L�����n��?����pBI��0ZX�N�s F1�5�({�hlQ|�D. ��ih_�ɯ�4����[Qm�7u�������zC(̗lm��MK���d�|Du!<b����������G5��_����d���(��U;Eݡ��!��FODf��`:�ۋ#~J�/qs?�|_���f�P�u�, �ڑ�Tn���Z�Z��1��s#����_��GY�	�� ���Jm����%���_�|�B��Z�麚+��$]D�p���m��	K�,�����.��m_3ѳر�j�ע�{Q��0�!�'��ͥz'],p�d��]Ep1���u�#�q�bG��-���gOa�4Z�箽m�>��c��vG'׃��~�z�hm��U_')�\��z�%b�}����Se�]<\-g;�9�4�w;�@�TQi_��>�$1Y���N�+��'�u�BA�f��ܪS!6�ys�\�!�J��Ţ!���{�h	�z	Z�A[�W-��W��W�Qv��LT4�~��握y��;a�o���΄�	_0�7�F����Z��O�׎���e  l��{6���D����H���m�q�͚	U�'�I��JV�:�-��GT"��*lx˭��;_���v݇?�W���y��D;��9�#|ޒ�`�M�9�#٪f��%-޲����S�Z�I-=V�U�|�Ç0bt�j�E�F8&ɣ��)'�� �r��������p����X���Q�V�a;��
f��{�ӣ���k���yjD����(.V�vcg��-*�����3 TP�5��p�H##X}��0�U@Ǥ|����X��ݥ����dL[���ה���Mq!���3vb�P���ؗ��:#��<���$��z5M�i�E���F�P&#AɆ�
p�[���ʲ���m�Vp��'.��lk��ߑ�gg�e�����edZe�VF�����7�Т-Yֶ��/��5�ua��s7$�c09�yo�W���q�R�����79�El3�x���`c؃�*��Ā I�M Mc�~M�?E��(2,�����&{�/w���=RG	�L��-4a8�K�,k&�7��{v��1�|����e�̎��a�{��mupሏO��&�s�9y�����H\�S&;����t<d�HT�*��(�=^v��"mf��s��3Ϫp�����.CV�&T
;���� .��(��ykq	h�������
���  m'Pt*$�˲���?(�!Hɚ�u_��+��,�f ]x< ��q$�5co�WiZ�_GM��o���	B�Ӱ�bI�"��f3����|0}�HY46���M~��H��H
SGRJ���V}���Y#�fZ��Ň�����'���/�1�s$�'a�UN<�Pi�_{T�ZXg�~Q�4N$���'D�C�]��0��FW%\�P��9w�����3�cN�ax��ci�u]�U������z(ݼs���F���<Б�r �џ�le1>Nx�#�	Oa�MS�[�;�"��OĈ���7l�?�sL� �8�̏�^6�Ah63��ڭl�da�)�b��d���Iڗ�@�#��_�0�ȟ��Ӝ�;]�߆!���LV��:OQSB��J�m �}-�_�6q�����T� R��I��󵋍BH3�G�ķ�5kEiņ�*�v�W�1&��R`8�\���<�`ߙ� ^�ц����✴A�Rus�v(@��ޚY�e��Ä<Y����� yݱ�ƒ���T�ο���S��(���3	����Yx��$�	"
��S�X.p�U�b�v�Y�4<�L�^WH��{�r��������}��H��!��黿[�#!�f7b�:	�)2��p�/�N�����9���bʆ�0Ϻ��5�PΑ{B��n������=݌�XD���=�^��sa/��Tf�:W��l�UO.�����U�M�L����qQ���C�#�[4�M��=,2a��b��z?8�V�V~�c�%�
�g-�8L�A�y�;�k#�|�`�(ۨ�S�h���C>q�u:N6ވa�z���\�U�����S9�+��/L�o�;]l��B��0�`#�O�C�מNB?�jU��^7)C/�6�O����17i>5.;O��^TK�IF�2�y�a���	}�|�y{�#p�g�!��#sj��E�8}��ߑ������x*ݢ&)�Z�~��1�;��6����J�������я<C#�p�vV��e�bMu�n_�'�N	!�jF�{���n;��S�x�k6���d����+�(H���L�=�0�4A͡x�s#����c'��:fVT���_�zS�4�m&��d��YB�!��C�<�/�K�0,Hr#d����pvM�`�#�YX�����X�@�"�:����{�|@�*,�W-O�����| �K%Y������4�.G�@+L����h��*8{xk���y�(�&`���UG��/G�����cGUXu����`����{�J�񌸇�Nv�7��L�� ��~X��)s7Vf[�F��d��k�Y�O��y���V(��:A�&�vF���jt��s�V21���ބػ;�krh� �aM�)���򇝭Գ썅Ȉ�V�n���n�O��T4c�C��7h��P+�[�b�\Ӆ[*�`#2c�ᙇ��y�k��z>�V.����}��
>b�1�����F��-��!@ܶ�n�ҹ=�#���';�s��x����5�m�7uЧu�R����cS^A�5�f;�i�Tl�DF�{���̰B���9ci6L��$6y�]��e���r���4��@Իf�'炫d[�4S��o��Gkh���ԙ�j����<���J�/]�C�v�щ�	�i��ZL~���,�/)F�I��#�Dr/[�V�v�*7
8�r�>�\,C�$��t7ņ� ��HX��2V��\�Xy�am$��@,�@i���4n)Fj&���nF�	6ސ`�Y��Mu������O${�s�U�t�QJ��F=�+%�r�Ď0],�RIӭ�}���#|�M"�1=]��8�%�u���%y�`���#L?��J\Ү 9�X�e�ǝq!��/oniN�s��庝C�W^���uH	k>���rV��^���Ax�GܵwL8��ܽ��p4a#;4�S��K���9Ԁ$�f��=@B���A�{��kM�qoS�i̛;�Z��#��cY���D���О#�]���34��旅A_��� F��D��om��+�a��\m��X�N��mV=@��k����������+h��)0J�Y<�)����è\u\ȹ�\�!A�_Ø��i�)�� ������K�{����E�q��Z(�Ӓ�sh�HC�b2ν�c+�ǧ�i���_�*%J����>��.ؚ<�ʗ��<	����*��)�)�=T�D��.\g��uS_��6F�_Kx��$.��<V!e1�p���+�/T������E���$���V���m}AƝ�\��fl���%Aj�֔H��qQM��@��� P�3�i����j�R=B���SK�j���8�nE��=�2�Sp���7�
*�#O��`g͍��_���[R�_G�'��E)��·5��Zby���4�40~��\��m.^ԇ��X��'��]�[rz�ׁ�lM'��Ѕ�`���yOf�)����*b|�q���!m�m���}[齑���(�ISW��^2����.l/]1�?�c�>j�����
>�¡w>2�ٚ����M�b"�F��p{6�R�7عl�t���0v��kC*�'���MRh'�o�&'AdAp|܃��I��,��Ϡ$+B\���b��@���/H��7�6��QF����HCZ-"���9%���T�b�u�rHߩ�+6�+�~�+N���N��u�3���3s5�A�Xc�K��>��}d�{���4|��!	�?�u�`գ6����z ���	CmCDfT�2H�"-����@RC� ��Q�|e��I����T��o���|uP.�|�a��]�7c5��u��,���z�T�;$MSe�rG��{�aB�GvE�xs�
�|�(�;Bj��M��-J���W
*�%�"s@�>�K����,�n]¿Gtg,�#,����&����Y�����:���^��kR&�I��_��;B�/jjhNcY���1-���(�m��Y����1t�����,E��Z�����S�v�ƅ�)����c��ߟ.ܳ;��Ǟ6�f��?����%O�w0��r<�tM�I���q�yAn��B��ꮧ$�~�'���V6�?c�T����Y o���*>OG��Q�79w��^�� ���j6����W`�öp�K��h���Ɣ%}7h�I���`t���}����4��,�LQtv�3=��B���(�$H����g�j�����@��J�2ۨ�
��ź���xW� �jل�i��N:�<�ވgۓ��#��<M�9��6��V��DUf���<���Qz��;�(��*#����Rd�g�~��x��HD�ǫ��͉�>肽��)'7[�o��nta���6"G����S�A>��nI���gߣt�s�"^�n���(�}|�����'~�2���`�و1����A7�j.iz7s�L2�Q�l��Q3zYt���\���1a����^I9o{��E\oɱ��O�%�8����x�<�*���'A��[�(�a�0�L|-�Jo�DOk�|:��2��όtqsYE��w���s�o�� u1g���^r���L0�V�|g�.���+R��}������ ~ѕ���A�7>���*�����Ei�S�#Y0ϊ�7%u:�-K)��<�|�#+$?���=먫�s�Сb:��w�r���� [�B��sj�?���nQg.�Ϳ�	^�a�鑒dD}2����s
�Uj���F8;9���h�T0�*�����o<���J��<�uK� i���6����G0NB���h9f��&�v?�m����I_����Ͱ��fԊ���v��q�_�YjS�k�TN���O�/�F6/�Q��_�$��aX�|����o��k,�ip�ӗK$�N�<�K��:7�r��E*H�I���ό�2Ez���g�����v�.��a0ϣ�яs����7�x���EV��tk�-��#���,a��aө�g֩<g��zX����xb�W�b����)L��u<��O��	_c���>5i��{� �,�U�a4�/�mI�3^�cީo����U�xf������A�
t������H7[؛��?�����+)��U+�hR�M���LV� /۾gלr2Kâ���ŉfqz֦o���d^�)�U�Twmd�/A�!"3T�O��h�&I��u�[�z�c8��E`�^����(�HV�A4������z��a� .�v�#�*��'_�%����f�0�� 3n�u��rENL��2���B-Q�E~]-�����l�
-d�2Glf�|V�	@@_�+�۷n�� -S0l;��_
d�̈g��S�c���:��#l+_��ˁU�E�������d~��T�
��]�>�>»r�~�x�m3��O�{st-]�\]#Nٽ� �s^N���+֖3xs<�tl��ed�:� (#5��5\&�|gޫV�G��xn���&rh:�1�ÆF�h9�}R�MXh����b1%`Wf�����W.j8�ȁU.�)ԅ\�rVG��O4��6�)bUl�]Y�R��1_b��b�鹁��ߙ&|�c�됥7���1Ё�Q����2��.jYt�t��!�Z4�`������� ���>��+�=}���o�t�L��F�^�����T��e��sl
�Ҟ��@��kc���4��W��$8o�!d�b�+�:G��jBJ�5N*���3���b2i�����.���m.��-�f��P�k&�}���8��}���O�s����7̮O\���=�(�0:!fN]���ॽ��O������"+.�Q�����L�]��}6c�ԋ8x����5R(��F\D#�LhKLmh�(ÿ�r�ڳ�B
Ш�u0G ɑ)NK��E�������n���ܚ�.,l"L�� ���������e�4�_s0;S�� "���8yO��5�)�X�~܃������P��3�w��|l��xH�.֍�d�0��|B{��D��JI*�p��M�~���Ry���e�dȽ(i�g�U�ș}�jх�_��`���&�*Mm����ђ�9d�Ho̷�9��5�e�3�]��ͼ��DJ��&#ĤQ�E;���M�v.�$��z�U���+�m��Oo�+;(�cp3��M�4����̕�*�xO�5����Y�|1��������>b�8��Cs!KSZ&���5_DYi0��k�i�"�g4�s�l�E����ݎ��i�;U�qQn�v�y�}Dה)!b��n�`%��93R��k���Dt���>�����I��c~s&���V��V=��3��ȭ���w39#ë��0؉���C����r�~�{%��6��-��D?��<�MR��C�Dy��kX��2�/V�oQ*�*�z�,���-�qXi��8DҤ�{�Ö��ym.� s!d���	^2t�PCMb�,ǵ���w�jQ��$}g�,�)�b��PH���񌃨���֓*��n�V:�!I�%�~\���4,��ЛEum�P7��6��!�q�ی.�1c��z9|TK�]�K�x���)�f