XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����M�+-㆚�̀�}=>ŏ4��`]��Yd�x8��'R�r=i�@B�ޚ~�b�_���X�ܹ�i`�}�[0Ǭ.UD�1$Z�k�8����K%ˢZ�5�Pfk$�FR��Q��*;(��@U}���P�yg����x�ؾ>Ħ̦���gt��#Fn���[��<
	�P������#n	O�F�-�鶪ˡ�+���R��o�-<�
��C�T�Q�$ �f��(������k�;����b߭��"'�kq.��h��ڕ��K%��Fɥ�6)Ě���C��)U�4C"�g�	2.�TH�5P���ӛ��v�v���<�ך�9ğBƐ�ɸ�����&���vxb�)�ţS�u/�'*~�/s�x���S���e����CH�:d9��}okl!�����m�@���iî�I�e�b��NZ��	����auK]�����8��ރĴ��v����I�T��AG��n�:M�8S�ih��&��l�v���Q���i�m�3�m�#kiZ+0�:�c~R�j\ѠXqs��3(���[�,�y0U�LaC>�A��'}i�z=��"�[Q�ț�+[���c�8���X�|Z-ʭq�F�}n�BtAlk������j?ҚF[攀�h���i������V�U}�(t�zk�����y�uO�Z�T��t�ìm�1�T�����S���s�H��
�gl�z<!��wx��6[b��(rP=I��D�Xj��̡XlxVHYEB    fa00    2d60ʩ��d�>�j��a���E�������-+|�m�-U|��t��l�Ӹ]Z�7�n��g}\0��~�T�}�&�=Co ��9?���3sH��(袶���� ��t+]�� ��S���[��M�7��6��~���a�Ëb��`����ٔyH�$�St������5xa+�ɧ��T1���0��n-�4f��Q�"�������"|�|x�>�s}�΋���2VqR�u��	�p�9�T�?�kݑ��I��¨�n� �b��4܅�g�L��Z���qx z0�0:ޣnwu�4��.�Mh�t�O f}��z�b{>.����a^��M}@8)ۨ�G�^�}��MD�)�I��W�vgU/�h���Q�Ҕа�Ѿ���v��ڙu���J�Xj�kP죯}�V&
�ˎ�
�g=��dR�zR�I!��Cv�fI@��*�?��tJ�J�"q�vI�2��Z�V�J]�d�����~�p�X�0�Ј�Cid ���	,��ej���N��~�ͷ"&���3�ERXq�BYj�7t�W�l��_pR-ⅫH3���)<,����[����.W[���H�D�L���ӊRW���\.�qa�U�x�|�7�9�S��vf	p������mh*;l��Mp�Br�����*+�j؜���^@9\c;4|���`�����)���e�m'�c��Kh���!2f�2[bt�*5'B�b# ���=���XћY������k��I����&)7�~+�q��W �rLl"�b�X�Q(Zx/<�I�{^�Zw�چa�8�y_r�����s�yn�yR�9q�4l��s�@�h,n��ʅ3Q3#�����p�� �Ŗg���!j.`n�\k�k���(KyS���O��i��)����T�����و�	gb�je�9�ŗ 9Z������c���w��^���e�D�Nǌ?����^v)Z_��:�����ٲ��E:^�Y@��Y���"3��5G��3�6�[P�vt�hV�ްꞝ������
.P�`����JCu�m��M�&�XD���,�	\4+m?OE���L��,�/nI,���TGz .Ӊu�t�b���onk���IC��u�G��{*m_iF\�}�V�	�e�;E �־�[,8�qHP] ����M��oؘs�F����]LG���[;���w��Q��f��t�4�(�@��K�L_#8ɉks p-���m}��q��8����>'��Lk{>��VN�7���J����Xp���@n�ٸ|Y}#�8>�l=�.ï�W���:jZz&�ɫ=id���
�5��5�	�f����>8>��A�w�D%��ZkW'&b����qӽt�8q�v������Z�D��k �<%�te�ĺ��n{x%�\ԓ��*�p(�_�E�ٮ@����$.·��.�[g2F'�%d�ZK�;<�����b&'�@r���y9�ګ�=�I�$���+�*�~O\c�p�̧�N�^�Q¨�m�5����Iyx�����e) �LID�j������`�*�/��,5�p*L1�{|�Խ{ѷrz���6�0C���hɕy��L[���͋��q%</e���!��ex �1��1*����]�{4O���L���F�{�mV��N���{�d����^޶~f\�mۖ*�A�\5r����z��s�"$k��4��;���9*f�]������#'X�&  �.�}�r�F�l
�
24�[�-ô��f�<�d�����G���y">����]�;��tir��FncL�R�N���,f ,��?���hQ%��GӨ�6�GZ����L}+b�i$��J��'1y���6�lÔA�cq)�X��*R�E����u�m���2�]�Q�[)�H�	 .�fs�VW��ap�h�]����7w<W�@KU+[�&�F�_b9"LnB�9jtE=
�S�Z��B$N�D��I��:mY!W���f��Ldp-@��$̶ۍ��J�a����@�g�`������o4����q�{9?�#
��;�@�ƥ��=eB�?�9)�-*�pJJv<?l��vZo��!4��e �+����B�?����*��t+,'Y�I�{
��!8p�wʝ);CVQ�j���a������4%V
m!�̛�rE��)��1+ΐ�6�MC�"!��(� � �tIs�̣��7��R�3EyV�{��cf@�28G���d��[I|I��lD%��
##�Ђ��Zf0���W#�x��1aK%��yВ8W]z�b�kt2�%�z����%�@H���K��a�3l=2��M%!�9����	���k"Y�+w����+c�@�m�6����W�v;�Ȼ �ߦ�����2�iw�.�1v�/�|��O���D�����z9\�Ĥ~�׆�qt����̑'4�,uw�ʭ�l���!'^�$U�h�D�(_�e�]��i��ӆ�LP�=e�N ���Fǭ�#Ax��N� �b��F��V�ߠ�Hv0�4���rP[QXwPG� 'E1]�$t3.�b�Q- ��>�_����G��+P�Wh����Jk;��ɋ�ؽ��y�޳ƀH �9s0�傮�W/l�n�p�'x1wBy��s{rZ��K*V�ƴ1�����\
�����Y*��K�?���$:���#��X
V�-��R�Bߏj�m���kE3��l*�?Hs��q¯X��.,��u��[l4��	5)$���V��.��=�k�Bt��&1t��=��	a�3C�9�>l��H�Lr��∃��o;�k	�$����iK����
�$���E�mن"��l�����T�,��-N�RC�݁�VΧ�	���R),��qe������絝��zv��)�G_ġH�P�|�]^�J�|��8��
��Ӳ��ٙ���D��}����M%��X����s�l:ؑe��N���Fb
B ��~��Ğ�j�^�,fbA�rމ�,v)F�A��v��@rNb�������󢮅:m�������Y���H��Η���g8�L�x$�w/��}).�[뛅��C7��Z�Kf��&~����H8�]��xC^�/yw�D�gq��3�_����2�R[3�1ψ>3�10��Z�W�!�nL�O��3��g�:��]�PL=��=����w�N{�c�O|�-@�7�&�]+�쎄�����j;fv����uӆy~�Wi�R�C<G�	��z��{����Ҥe���Fb-���bU������V�����k�T�>�<����rJ��g�?����H{U�+_�1,���G�l���r���AN�F�A��֓��7H�����(�\�~yC���C�;L�lel��~/*	�P/nE�+�a�=�E)�ؾ�]8��9�K�2�;y)�Q͔�l��!����F;�tjO�3Du�˒������8[�Q���<�*�qo_�|J`���g\�D(�{&Wj�6��6zP"��h�;������֓r������x8��m���n	�W��E�F�h�7ذ��f��j�z�VT�p���6��L����h��V��e�=Vu��.Er�qx��s������*�^/�t�I�,�簵^��"�j�S��<v�Zqpg��J�-� CMC3�����8-���y�K�I��(�HK�h���(/>�����]�B�QV���u'��]}e"�5�������t�5�J�R�wE�8��z
p�a�ao�� ���Ǭ�R	��PP�o�>a�I�`�(=�΁21����R�ZC
��������l\���Xأ�T�tu�M�=�B�ǧ0wv�M�V8H�cD����ԽiW��Ӱ���P�zr���T�1C�J���h������Y�� ;��d/&e^��`��J�����RI��\�N-��,d���? �ޡ-��<�cޢ��)7�E�J�8����[ki�z*d���U�ק��t�}��j(V}��w�#����w��mPB�pk�'U���=C��$X�4s0.X�v!V�/nF����5aO�҉��՚�mh[��t�!��`ƪ��r�d���W�O3D.���WC����:�4$�X�v���Q�*+�kvs�CK���~���8��+�|������UWMj/xQ�Y��SX�Z6U&�N���|���=��p��.������o�A�1�IKn�z��U3ݛB��4v	�4ݚA^���š�rg��� ���Q���L������Ѐ�@k�^rK���[����#�M�>;�zyNrs�a;�E�H:^�D�F�\;Z#Q�6�7�s+K�z�PK������}Ǜ�Tk�}�p�{l��ɬ����L�3�E��B:Dh�1�� �T�Kҗ�Y�>��og���EQ0dP�W����<�m\�)��ēo�ͮGX��M��;�m��[�,�E�;�	$�P
HSF�܂ق29�����'��wC����w�����g̘�N*�m��~쓄^wY/��5,������~1du;WH\\ �0�\b2'��O�Kk��*
~2�,�o;�$+�6j-?�%�q���0�lo2���8/��"��/M����vE���Ų���*b
gX[��@+<���[�C�
(M�X�+�/_z�ۿ}��[
27��uf����>�B�D��o s��� ����ֿb����a�6e�;D�8Q�Y�^��!�y�Pn�1;��y�L!�s'v���)�̭{ds����6
����t��x�E��=�F+�aT&�D0���|�,S�� 4��!��U���	~�F2R?�Q,�-��t�X��'���YB����tP�I�瓍&?6��K#��+�(��%p~L�����7R�O<U���!`l�W�]��H���,��g�#��}��o�v�m)H�;��驽q�qxn)F"�������������	�S�G���>K�7��t?�����K�zZ@"�:T�d՝.(�g���ƅ��V?u��J!�&�
�����D7M�q�AoP�J]E[��̂S���A(�&��y�8x�W�����E�88o��f�N&�t}ɠ����;gň�ܨ���Vi���0(g� Pz�����_s�?����Hv�����q�+)���Nb��"̣� ��pY�����N"�Ǜ����"�_C����'�J4	F��A��2�l�mQ��x���ZL�4���5/��ƣ@�t�`����LEPV(|xn��K(��qnb
>ʭ�����^���*����S��O<�),2����¡�9�d��\�Gc7���]�S�	��yi������ف��P3�~�Dl�E��z�`�ӣY�1'�=�I�=-�\��O/y�H>W��\��8��+aWWs���X]Ί��dv��7Gq����W�=���rD@��Oh`޳�8��r���茟;/��$z�/�:����v����KQ��('��᥍��5��A]$6#`��	��<���z`f}}fI�#�`�w��>X΋�F4U�K~���M[�:M�P���	��d:��msٶϲ}�����*�T�? 'T����W���H�%�$ @Ԩh/חۦƼ�/���[���I�V�i�B{�U�;#����Gɚ��W��`8}(�����`���������ƪ���uஞ궉��-����Oy���K[\@���� ��Ŷ�f"�3���G���3�I���� �>R�y��c"X��>){~Gj��_9��GE���k���{&�%����Hp�B��y�j���@��6�T�FN���|BRl\1���W�l�lHGg,��ER}���![V�tT�1���^5%J��K��s �#4���<���01g��-6o�W�L�`N�Y��ٮ��8$��S×�̠�ζf=9�:5�ed�jz�Unb���H����I�`�ّkD�@�I��]i��,!oF�z��}��v�do�����Ō8RH-b�/��o�ٕ�]�G����M^ބ��:����`�O$s�_  ���Q���1ѐ��cnl~�va#���_vӨW�=bC$^�v�u{E8��˅(,��(��2Zz�-u��%��bߪ���o��8�M����ØA��i�!ݣ�SN���*�i�eq1�K����|?ej���qW�͹Z�bc����;������*��1E���Ջ�q�O�e~��b�R�ڷʤ$�s�x� r .���E���j1�+.�v��$��y��KA}�'����6��552��b���J����D�s�ey��`�X�%<�H�+x��z���έ.q���{��{����z^�4�<��@�$\7��O���(��Y���X]�J��'Q$#��y��G�ok��A~���:_���]�F����י|�A���4���X�ar�n�3�ߴWFE�fw�h�ڛ4����WZ!G���K�&���D���%3�ɉ@5��tI*��7,����/���[93f���hl^Z-�Z����ޅPlpK���`���3�h���ĺ)��+ݑ��Ⴊ��$�3�~��ͨ�ةBWp�s���t���4���=#+9�7 u��ی�6) �*�쪉�k;u	�}*��yڗ�����o��G3i�e�mB��-�W����Ӣ1 WN�a�{�p�Fc��'m����y��z$�����(4(�#=�� c#N��?�V����s���0�?E��r�`�Gʟ���8(��k,������#�\.D8�d���]��L��{4g4�f9�pZ�ɹ%~&W�����vu�]\3j�7�&-�2�Ƶ�=�L��l�>?)¨�`�Fh`#z���%ܷ�ʃ���ꨬ^��#��SuJ5c9�lN���L��H� 5[C��u��+9f�Ⰺ�:��:�7��.�ꥌ�/��ei) ߬7�d'�,9���ծ�⟇���*���J���e���o�k��ĤŨΡ���s[q�]���)�,k�D(��{�q~[���ȻEg��]�
�2n���b����U+ڃg��m��LG��f��C6��Hf�U\��ET6������sބB*c�M����*d�hQ+wa���F<4:�s�/��}�fό�#�kg#}�p�����
����W���p��g5}Hd*�Q8̊�y���b"�8}�?��pp�U.h�\K�wmO��5�׌h�eC�B�6VR��;��U�ϲO�J�U�? ʫ�C(,�]�"*s�2�� ��VV-�Y��2m��I�_NEf-�	,�Ƅ��>mU�B<�h����N���+R��!�;p���w���l���I�S�^aCĩR�	ݵ�,���D�=O��s�D�w@�E��Q���+zd�*&�b�
�n�{�1���(A� -������,�'d�Q���<��l�:��@�2^����3(�	�Y�;���*mi��_Ú$(�_�K������V`%ѣ$�M#V��)���cP<�MI6����#��H�T*�4�1!tw������#�����TM��W����
�5H�h�:zV��A�w��Q,�h�g1����-.�ō�`�$�*�6�	���X,C�qi��ꋍ��?l��1n{[<;��Ͽ���hY.O���\�6g�4�ɀ�gh�tZ�OY��{��k����幱ww�8,J���8yf���WDc�d�7����������Z3g�.����j>yI	<9U��)��J ئZ��2d�wG��s�x[�q�����{�Iٴ�Z
���a�������w~��,���-����
���|�PpED-_̞�.3p����}Բ��?x���~;-m/Us>�x?���zf��+�^[�۷/^����7�����U�9�M�\�M������ܨ�h�N�CѰ	�F�y��Ǔ�(E�zuv��~F��;��Ín�i�df�22U�ela➥���qSs��ʚ>�Ǽ�� S�����IMk��K>��`2]_}Ou����Y���ҫ$0Tzh�3v�Bҵ�U��?<�i3�����2���D��	T�D�^	 �}!���e^��Pˑ��7���6��W&Qӆ�>'LꅬsT����_%����NV��~·�{������DJ���S�%�tۧ�35�,�$~M�,	����~O,����/�!�!�D���2>�>1�U밣���X���B��Nq�$l�'�ÔFh��:k�����2����S�Q��ҋX�W~���r:��=��ݻ�,|�cSU�"�,w�qX���~43{X�6�.uI�QѦ�H���x���2��F�7�O��N��z�S���W�����~֐�l���P�&K��L ��]+�]�D�@iގB����*Ks�*[�]��<��r����D��¯[]@7�>I��.�����d����X�iuPDg5�����l��t���67ح~i}�s�1�A��4�ߣ5>��?f�"w�|^u"72� (ARcǱ{a�!�_�Oԣ�#)�����A��dT�:!�nm	��C�g�r���Ə�r�)�0�+C)a~�D���]�Y)����x@e�܏*x>7����y���#c��(��엍��(����A�Q7��&��-qmH�x��G;�LK� �T���/?����^ֱ*^\�XG
��M�z�@�@l6B5w^��]��Z`� ��EMQ�ޢ7�̫ʫ�M�f�s˲�H��Z�'��`��hr%GU3�����0nD�2���m��|���(��P
*��3���nn�u7�Ii2U������z^�ƘF��g�G6"K��vX(D�|d�����Cs��>n�ch(
���	�������'^��p�5!��P�L	����j��.Ⱏ*7���?	A�����#*�g�����a>xku0�Dx�DX�-��Wo�ޢ)p�>�J�X�W5'��kȵΘ��C�7�D^��O
�h���3t*;�������y��r෗��ve�P�Hb��N�%6�EE�5��_g;���˙����6�-�?������������_���p���2J(U�~�e�Т��6�O���:�u2)WG��e����5`VӲ0ie\tQ�͚��{��x/��0�8�VDB�0�m�������)�����d.�-���l��u�:)M��M7�Ef������s���f!B��x�K�3�'M��I�XNbO9�!������u����Ө#ICA�%Ȏ̰
�A�o�N�����u�������x�p'��RuHH�d����;�.��bD6�n�;gC�q}�� ��{%a��T����!�+p����Z�>D�]\�P@�����a�tzڰ����$�;6j�+߯�ߑ,��ŗrF3�(�NS<�J��.�l�L{���@%����3��4�t	ɺM��#t�1�Շ�M�B@��Y���v!Q@ؓu��ip�k'j�vd=��+�9}���I����K�܂2F?�
�n�u��P-��ed���C���h�w׀gH�"��Ձ�H"����篔t8׽b��OU���rX˨;�|�D�,:��_:��M���ಝaG¹{pp�	�E#��#5��|Uiha�R1��t�~�>�u����_.!M�0EY�ju(z�tĻ�L��<� �pXŎ*�SF`�dWYn�:�sg	AM��#CB�5�D��ioO��|޴�qG�s=�܅��+,0���
@&A5�;k@��b���ě6�����Pp��lW�03|���{D��PH�8�v�;�"�Fv��F(
!i�\CŁ�tq�N�ni���3DW���r�Z	��AY<z���V�1Un<Y�L�7a=;�x���)� �W��Mc�p�y6�适���M�d��\�F�
з��}�����h=W��T|9���>���4�I�FU:���ԓP���99j���3������q�h�S����^d�Q�����u�@�f���Z(~�L�a�a<�+2"�t]��#�?~$�d�.ꅎ�k5�8��՘j+�D^	M����*��M�����M�j�s5���.M��<I�(0�K���N�\.��\=h|	�E&y��S��t���eW*��oC�0*�jSͯ{=��I��4:�p����k�'z?���Lk������͙w���C��%�x�����T!}�?��n�k�5fO�:"4�S���k���<���������j<�F^uhS�ݬ�ճ�ʴ����b�j��u*�Vxf��������1£/Aa1EP�����vI��[R>o�(1��PwN�����|���k8^$�����^[ ��q��@(���^F��ng%Q�O����C��7C��aq~F��/T\.g��)��.g��Wė� J�6V�B�׳7w0��!wp�W�+F�5��k)毽m�lߑ��G�TH�~�Ift%:_��q��i��d
��V��Z��yw����(��ږ
���gN��+� &=�"�RkUh��g����Cg��z c�D�IS��M��DȨt�j�x���:�I`�X��:q�w��\I��Yl�akc^��y;��4�������)�D�����㗫���E��b��=,���G*i�W�uLCKк�9�=�Q��\P�0���i�k3���e��)C�'��K���؛����0�HC���J���y�(�pGc&�}�̸y���mko��
�='�U�֠\�6���y����v�E�����s��RJ�Sĳ(Ի��J��/��gӳ��\I��4�"���`�1�=o�6�<�D����s���?ge�\E�*^bV�`U�8����c���:�����c�5�0e~t��S�(3|�l�]���٧�,���T֠�z�N�pNH$�!���$B�IڣA�l�U2���s��Vr��N�NL���D���P#�Ś��B�����~�W;_�ifơE�؝*�+�ʆ�l��Qǡ=�3U�\��@l��� �ϱ�-u龽����F�A/�δ"�&���c 9��ʐ��Zޜ3t�,�Q��Ճ`'Ye����j��Û~��گN4�33��:-���Rt�j�4;&&X�Q�vZh=lYQs0���.Yr9�ú�0�����̼��&����oRՔ��%艁�t��tS�l
���~�%y���ה>P{����BHa0�j�̾b9-�~a�<���b�Q�c]�\����l/�L8��b��I����w8K�J��S�C�!e�L~L��8-I�?T������s�ĥ�=���K�ښ�#�u��9��H����F�/�4�\�+�H%����n{(5/�fg��@+X&��7%h/���99�Y>��
C�Ԁ���Z��z;���E�0�q�e�Ι�8)
f�7�Z�߇0�8�\�g�9v�(�h8�`�fL�4@ ̖~̓�:�m��]^�IZ2�uݞ]4�k�������id�n�`�F�
+I��XNx�~kO��Z��^8������@�	=B��*ax���=�G�?�v���0nu��?S��/bcq׹k�b��A��v,�d@1��o�-;������+�lph�S�)S� ��!y)�K|��XlxVHYEB    5914     f20�D�z�1r������}.�UO��f����T?�1��8��k���m.�;��Y�8���%e��g��ƥb�>�!��N+�xƂ�����S�_f�Sl��sJ\�"Sd����6f�2㐭���~��;A���4�u�q^ں�jK����I�H�������awZ��:Bz���.}�[�AĊ|��{Q�4A_,�s,s^��0^��x��cbc�*�@�S�0؎�4Gf�=�:�I<��g6�~�q�3�]\�p��q�"#�D�#x��h�zAr�6H�sOEʡC��ǹ
^ +���b f(I�Yo����w�"���:��Ȏ��0A��q�2{r���J���DY�OFq���А)(��΀2���/�,%ڵ�`u���>Gp{C�6�jZ��ɒ$���A,�rn=��(�V��	� ������ѯ=��q㏔ �'��ml
i�3U؃L�<l�귒��8�m��E��Vo/�-!�(+���n⟲��� �.ɧ�d������k���yݨ̞ܝt�lnǔ��$âjF���C��a�m�����4�"r�b�Jk!3��kW��۱N�_~�e��u�8P�|�Ç��X�t[%P���r=�7�<� v�f^߽����Yj��Q�W�����W����"t����� \�A���$���8|;yT^���������<��s�� �k�R��j���`���\�\��9��ydQ���/a����qB�~F�b�NDH��C�s�&ZZd5�b���!����)���m��ѕ��Qj+9��>��Ӯ^@K�6���� ��~�/ڀ��~�w��蟥�\|j��2P�
f{¨��x���ۨ� ���:�׌�N-�A��I��:@���,[5���!uG��|(�(�|�S�h6u�+�RM����ݞ�MxT�9�8Ʃ�v�`����D��	S�_��k��w.3:)����?��c��)U*�A�G�������x��y����J��c�U��&�({��8M
�E�Ko�~�V����#�����4P�| �dX\&l0�i�B�,�+b8��&���f��)� 
}��$j�~2�����B�LB����L1>��[*�hN�2�Bb��?���aY���= �B�����`!�i/V�%�K���i���-D��yzN֛ht�T����R�^O3�	�g�S'���꧍��C��sΨ���&�$��y�=F�۝KkvkkdŢ�v$�WS�����/=��-��߉�z�|L�#���)����DA�%g0^/�dD2El�⺍�Ǟ�"7�u�X��Z7��B�lb���9mZ�A�y1;�ܩ����jsL۩Ȏ;'��5z�B�s���rW/��`�h86�b4yU"»�B-VP̳G���C\����J��!��`i�n}3��-1)�,���,�㞊G��N���cO��� w�0NJ�	kZ^������)#����!��p���QذI�������y�b��6+7�*�2��]P�J��ت,5�a�k�� ���GE��/橙���C�R��ʄ�60�Zܥ YR��Wv3���1ME�2���2/$"2�&����MA<�ZH.�F"�o����>��楘�Aj)�G6�{$"g�y�z쌹ʫ6[��W!�PB~sGE���Y^Aa9�[��5�K]b��x�u,�f��9����Ui�(=xvh���N�i��l�j{y4���<M��WY�c&�'Ң#���x�'�M�`�e����q���|r:���t��9�Q,g����PE���S���e�N�!Ɣ+Ћr0�VO���*�aĵ�Z̺{�>Oh�H��͇-���B�=�	�ￄ��ᓒ��/])o/��ۓS�����C�����)F������8�>���k�и���K�=�9[�Y�%6����l�=~>��ۥ�4�G�I�Ys/v��4	ؒ��y��2���@��ϖ�i�wޤ�ڀ��e�sT� z���eʵhP�ֈ~b%*��u��$�#�:j3�^֏"]T��͵ �P�x�I��b>T��0ܪ;���S%H�=.a��pQ�#�D���TLDz�]L��)'�;:IC�
I�U�/���D�*9���`"��4����z�l\��+ˏ�v}������:��d}K��6o�\�TР����Uw:��+�:��!u�l(��X==�} <�T	8���_��Ir5SU��SU�B�
繆�L������В��@�qB�城K����X�;R��VX���	��ab5�C�&�� ɵ�T����&��1�3����z��b�,h���L�v˧敁RL���4�*K���N�F����k��ӭZ'�u�V���ʍФS{�v��F\���qA3i	H�l9�孇M;�CH���^�E!9����l:�E�ٝ�b���"ӛ`�g���k�_�� ����1� �l\~
��|�N��]Y�l�fƶ@�QL9���S�����a`Z�~7[C��taUfѴ�T_K#\r�f�b��l���q|qY��XY�O���]9:����%�i�y�����f��u�0�Ӧ��)�kЈ��<�)��xӛ�cF	�GlVB���`F����`��eɪU��3�H�V���%����D�TsR�,f25 ������`���!p�p.�MW�-��P�8:�lΔ��"h{\#7�k<LR�wp�@��8�3�3(����6�v5��h�٢"SId{DX�JVO��J���opI;�o��(�� ��Na��YdYm�����K�����4�ȁ����>,��Y！֨���J��Ƃ(S�/���%v��Ҷ�b�(�\v&cJO�De3�J��E�zNk^v54��4����6J0�v	l���LVgg�V����B@�j�k"�-�����*�ve�6��	^C��U֙�*J��^�pҿ�fPU���g	�jn�Ҕ�+��'<K&��������Ƃ���?/Rn.F��т�S;6M8.Ntp��pv���e�K�i���d6;1�YC��{��Oϲv��f/���Ё�x�v3ʌ֍�g�0Q�|Xc��Tw}���Pȫ����jUE��sw>�c�3�[xb�%"��mԧ�ڵ<[H�
3mx�� ܄K!�`67"?m_��t�Ս釱�߽y���U�Qa8O� ��ྷ)���aܨ�=E���1k
n����]�FD�0��J��.����-�������Z���2�JiU�ׁf��g-"Ѥޚ�i�����W��;W�F�)���J��ڼp�-`T�(�66BһZ���B�֘���d�=R��/Z���l {��@<�|�I�Y'`���1����;\?��T˄����Zm���U�Z��
1M��T��3_�!�.�r��NHYQ �uS�d�����ZkJHV���Jy��I�]��z�'��t��5C~,te��h$y����3g=�{����d���Y�Q�$+�0^�7"���J�ߨ'�\�d
��� c�g�D���.w���_��45-E�kA������j��:�.C�Y�N٩�D��Ϣ�' �ir����8'�B$-��_
�+FOB#bˏ��Ґ��j�ٯݟ���1��qg̾R���N �&�t-����K�������+]�����I[
p<���~Z�r�����m�NIb�LĨqQz��%�&����	g�w6�&���vp��`3�6+�N�a�A��.��{!k����^��uC�9}r�/� ,�f��X�C��?c��nfZ���U��x�ɵ2(H�?�7�c�B�5w,�Qk4Z�{�Z4
�֋@��<霦Դ��\��[���읰�B�<�o�=U��j��aEA�Hb��