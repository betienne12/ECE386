XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�7G�	B��]��(��%+�~'��>�{��2��>��(z�>�x&��I�.R&g9���LW2�o�W�mӠ�� �p��u�v�����_�_�Q	B>�L���n��ӭ�@8MB��V	�(TV��}4�E~X&��3<�q��U�
��K��Y3��Rf��8wA�J4(P��A
;�6`��ʧy�G\�N�`5��I�]d/��XJ&&��|��|c�w�EϏ���V�-s>i���wD���[׼�أI��p�Opݸ9<�p+��|���w,�Q4�i���ub҅���m�F��(���I��Fg�zu�c�Y�OS�r|]v� �*��"��ҵ��Y�ʥ/I,�4��9��)�fr�.(�ğl9'�P����'��ՠM1���i��H��T��.����u�uy����g�C��/S�y���tU�c�A�N��V$Ӱ�l��߮��[G�-�w����f��	�Z8L��FL��01���r��&�{���6a�dtᗀ$���vr����Q˱���l�z���U� ��դ�Yf�j��o���P���0����$�N5��4ߚ���6q�aA�M��rF�F}��q��F�w��<�(Nq���8������II���؛��#G��j��{Q�u.�s���W�q��mq
P�tK��E�H4���]R��L1Џ��<{� K�!�?씻3�������w�F�����L߷:Z'?	4��iM7�1"iq��XlxVHYEB    fa00    1790ͧjBs{�v"!�A����)�(o� �MO� 3K�o�1L��<-#b`\+ΑpZ㗲�FX}�'���M���2%��}A$ �[�jEs���swS <Z^�/��G���%�!Z!s���4\�>H��Yy�1ݐ�r�!w�l�H���3�R�~bR7��ռ���a��W������=Υ]cIvPk�d�S�O�uL��e9�8��ͤ��/��&,S�Y����i��5�&xX=u���k$V�;�DwίxN��3�����TZ�v�W૜N���8���,�DZJX���&�ǜ������q�Zi��W�P�>Z�! �l�6V�_��GF� N���T��r�ss���&��R-�G|$�*�V�Q>�C�dq ���W~F`㤳Ks �C�QLt�'�IŤc.�"�M�qj���5�r�Ŗy�<��w�R�I�h��+*p������1:���R�� ���L0�X�L���y�N����,�]�P��q!�v~2�j�͐�k�=,�>�lZyz��'J*�s2p�`�(��r9���rua�;�@Ew���K�W{���76]��=( �
=)
�O��[�zZ��?g�,�c�&�zj��	Uz��Q���qg)�
�f��Ϯ<�v���8bhF��ӡ������f5���0��b�Y����/�F ���B9���g���m��e��[I�1Xj��V#��KZISf
棌��f���/b�j ��pٶ�I��*P]�!	��/��=�� k�`�jF�1�����a0F~)Sk��x?�.=�6�`��L9om"ٰ����0�h��H-%|�2�������Q�G�I��[
̂9����n|m�l��9����Nf4��l�Q�rH���X�<�� ��u���,w;�ZX�\�9PJ,���(�5tK3.�8m'�̼hq#~U,u�U7��.���m� ��:����]:�Fc*��R>�i5[B�0���&�n(>������؎A���ݯ��ek���5�z�p�4Wv��>�G�w�u]�Z`��,���`�w
e��K�9������Q^���21V

t�2ĵ����>��������WK��v�0]Q\�a��#m󁐶�`���� 3��
R�(D��������.G�v�s���B���p��x�Xz
�:	���ߊ�����G�P<���]ܧN��� ��|,:�z^�Q�@�+�R��(A�t_��t�Jk l,��J���N<�g����D�Sv�%ޔ�Z�5~���}x,�r�[�
N%;���,4|r�G0.��.����~fE�:�.U6&�H�9�,<)$
�������G2D9�zAO^���:����%�M�M��Q,��%��w  -���K����3���^�lQgp�Lp��)4�r�+�E�^p�����	���=3��������p&F9�ؔ�1����G�O��;��W���91�x'`b[�_��?V��#Q�l��P+�'�z��ŧ�umۿ(?ݘ�R��m2�[���Z{��7��)�H���PM��~+�q7"[ﲧ�^�>���F�z��;�C�,��@E}_�!;pi{�ro��JO�(�9RN��,�k $`����;���Vl�h��|���Rw� EH1�nyM�-X@��v���^wÛ����W�y������3�A^5Ld��\��~�lA��A����a�=����@��a�h�R��*Z[�4m-1|͎l�l`��P��؊
�5�c�.��i��6���׮�e7����/D��a�P6�M$��9����?����/��%�j��	�4�'B	:5���S�hR"�/�˺p�z�#L��1cKX��<�b�GW� #�"%����Q���D�3�;9PI�������J�C��hr�vi������,ps'o��H ���l���A��#t��&3׍�KA���1�j���nx�Y1b����c�~�CFB)�W�}����EF��FJV	���ޛ����7g�)0�HA �x�*�mb66GU�o��P�O��<jZ},Λ�Nz鯈i�J�
�*5�/���F�<�@(N���	�t�!����Og)O?���@b�w�|dg+M��ᦏR��}�8Г�/K��i�[�\^��n,rL_��������J]��$J��g�֊Yx}�T��nb����T +*=����\M�,�b�;���O(��Ч��y�m�÷>g�`!�1Syx�u�g��TKXD�G�Ks���!A�`x�mW�qFr>������2ul�痥="���Ե������S�Ex�����3fc�����c	2K��ɛ�i���Lt��;s����TP�{�����񩵻��(4�zy߷��"W�9�۠�P���V��3FՠP��z(�|szS䯱@L�5�x@��X�
m�*=CD�Sk���z��Y�L~9��V�v};�o#����n�20s�Q��~(�Ӝ�x��w��K�T�N^ޤ�Ԥ�ͯp�!�L��.��S���1l�kL�Y.��3�(�>]YysoݨczӔN��"�����en2����>��^/��	�"]�$>��}��Y#�	\�s���G���8���m�Y��/�uK��HN��h"�tF����E�.�_�m&��8Xb�"vj�U����d��颿����Dxr�����.��qm��~�&�A���BS���:
��Q�pŉYvH�_�x6��u>�P�FL��$,]����b���@w��|-s�=��[��l˞K�OP��u����j�y��W�,�yj���l���o��pvL(��ǄFf8��{�?����3��B���-��]�O47] t�|����ю���A���߱���a�6KD��E��J�hQ�#�-�Ƚftކ
$R� ��2�q��0������.��Ŗ����v��dթWw��G���zު��-U��<�.���f��uWG��0i��P��h �z����S��0q=�����,|f��������4�B0*1:�
4ZiQ��� Նl4_�/�)(���υ���1^k~!/��M7�9�~�8����O���g���4OM=���Z�)k��0�K��� u�p��+Y!��L aT��Ə_�YT�}vI��/�������i=�'c�2?g�+�7I���K.� p��)�QK~+��d�b������
�OV������C��r���WX�B�ĩ�|�f0k�tH0�	�{�0S���2c_;�m�m��!\YEc�{ؘ��]���q��iJ�nV#O� �75>ZfI^�<�{���	�WqߎBu�Y�EX$N��;�J龨p��W��g��-=��&x��m��qT

I��[�~�xP'Ԩ��f����?�'��U�tp���+�p�=�á\��Y�I�\���[�@�J\�~z� �ŏ�MtrҼ��W*0r�G#\������t�O0�#���L�M��Qc����znw-=�TZ:���Bp�%��d�=0�'��u"x"rYm���L���%#1Q���w����ٰ�����ˏ6���9�W+t������E�礚@�fr��}o���A��:E��4�����BDI�Z��}�&��c�(n�-K���":$�9�)���,���*�n��2�Q��Jt�D0P����!o8�6��5'�N¡�Մ G�$�)qQ�^�R�[v܆F��ހ�}�J�Zy�08v6꤅�e��́s�B��.���V���B`�u3	�l#�L�ɟ��Px�	��,�i��)�>�o�.��~�v�Bo��TDD��A����ƻR�Rg�ު_�3�����A�^��ER�*��pxɉ����a]�Z[.(���^�V{z�JU��j� ����R87�K����	B�.��ȝgF�
|��m%ʯ9=��z��;���'�ZD�uǌ9�b4�?'����5�J ��1��"�g3��[ym�q�����U{q�o��98�Jh][�#IK3�� RNѫ�l��`�Sb$� � $?����f��Jd�UH��g�S���?	p�Q�w��jU� q����� .��b�D,��WFy���%�s-�{�EC0�*��X����M�T�v]��`����3;����;OG��f#䌣�
�q����]�
Q��#�=�9�I���ڼo��P��LF���籖�%��F��r�����A*�r��LJ�C�?�?���>�t���ypUrW����
�4J.�n"a�!��0��� Ռx��y���G�����a��!K�p�fD�cKG�	<��9��ǒ��F%|Q����E��!.>5otvZ&�ň�/U�[�\R��p����"�T��<Ln?�؇Qݐ�RGxͬ=�5��C��y��uW aFU��(�,��x{�Ǩ���5�i�����ϻN������z�5g���I"j�����˫���"S�/��/�p�	±͐~V���6��(&�dc(���eL �@ r��_13��gr�18�KҔBljRx"8_��_D`"k>&��e�IЃݿ3h�9�� �`��/Q�h�N�P�ӑ��S��`�[�%5�ܚ���rP���6-��)�L�$QֈeMo
w�Vk�����b,�\D�t�,�z�ԯK�G/%��'��|�����᤾'�6�Ӈww�I�'��,�q*���W$�w)�L����n��qu�Mu��[n"�)�x��HӈO���+�ٶ���?���O���p�ye?�7\��Fv��ms/�,���B�D��r`Ŵ�۞����ů�>Ղ(�����[(���t�b���E��A$�e*/Y=�2�p��8Ga灧v�@çf�C�����fiV�&�U0��"��W�p�����?V���U���."�櫔�n`4ᵟvwV5|6 Mi>�a��׮�r�H���_׎�{��P ��8�	zv��X��a���My$%�	ɉ����D�D��.{�F�����H��O�d<fQ�2=��oa'w�!#
�va.)
y�*}V���uk�H�����6�_BeM#Ss\�)�<��)0x�NvP��6��G1=�DOm]JY3p�7��e��Mᑷ�+�i��7�
RK����r�/Hԝ'z;�9��

�Idm��"�����6:w1ΗJ��Sk����_c�n�=����5Z�
���>�r��Ĩ4���<�l�>c|Z	�a�ˡ�J��Rژx?ډ�׌wQ攕/|D��Z\�3���0�O]g���Hv�-x�6�5-����7i
�-�Mb1�
*-���ڐ��5k�_�j��V��Uc��}���d��z�vl����Z{��R̓Ryz���Q��:�w�-n�ua�g*Rt�r贡���j�O{7>ղ@4!�A�����O+�Ŗ�!
��</h��8�;�����~����C���^l���j��N�	��Ѓh��M�E����RtZ��@_�H��HǶ��Udu(R�M�z��c2�D�B>�$���F�c��e��J,n���S��y�
�c����OaQ����2�~\P=]�2��:2�/��T\��>n���|�d��ka�SL�(O�0�+�;�q�5��35_�A_$}���/�m�4�\`Xob@@�������<Vv�8(f� *ʑ�i��p���Rq�{�Y�`L\픸L�՞���ly)�����,Y��Aq#O~bǴ�J�����Z��<8�/js�9K��Hup�D�X��s�Tc���S_e��M:�+k����z �@�:�]ē�.��{v&�E["W��3O} ��~�/~){x�ܱ�m&�v�N�~��>�t̂���y��K��^x5��y|�i�a�Y	y$?��Z�"5V� ���_x��R�~���2����m��p꣚V�!��� ��EC|�:�$���񀓨���.��{@{T���ztե�+Ǔ����bc��QSLF`XlxVHYEB    fa00     5d0;ϧKƠ������M| �����D�}�U'g�E���M���:k/M�/G|�:]�t%O`�%�X�����/օS$�w_AR�{�����l��^��情��DBFt@�='�����[��y<��Vn�BSH.4��F5o�I�K�2�^���r�za:@~�����KX�~��R��0�K�x�v����Q���\;��8��[�=[�\M�\�dh��E[�� �
x\�k�$�IU�u-6\@��"S<�ELTXlP�&'���S���ml���,_�P�ԉ73v��y�N!��R��h� }�쭳�Q	������M��CMHZ�($"��+&U��ʓ�/j5C!o�?�Dn<֥�T��V�??>�pVxT�-��-'a�O��R���H�+��B�����0�A#�q~�2�����7��~�+�<Q<��A�b�������!��Ρ�s{S��H)��Z�M��N�8�u=mo��+�����/��c5�{�%���ҙ�k� uq��F���r�kL����OV���7~Cz-��8�4v��d0=wm��!Ґ.l��;U��KZ���Z�=r�[�f>d�s���CUp��k<�9�s�Ŷpc���X�ᑌ�H`�����������jҲ�>W/���ӋTN�0���#����w��񃊥YR�|�n\���Rxxb��g�(�V=�̳�l��j�t)���ț��gVi��:�A��}�uA+�e�:���L '�,\D=̭��76t��S)�ðS�e8���g��J�������4a�������A^���G���0�5�Vp&��J�2�TdQ햳5� ��h��{���H�ح*����� �R��Z�k��ԭGS�[���S��\܎j��E�iYي�>�e��~�ڵJ�`G9�D1c<��RC�sj&���QIK���m݌qH�ǜ���)�Xہ`��$�SI�+�ERڡ�}lXX=�N��|�o��Q�c�\(��sß����{		k�kWŮ�ט(�v�I4��@)�$�K��_�6!���S��r=�����c`dvܗZ�������D���\��Q�#�h�E&@��;�=;p�5U�݀�]�i<]c�Fk��xѰ��F���n�c�l:��Q3�����ީ`j�
�ozFl2��$�G`�IyT�f���� ��O��C��Z1����<)*�he9<T����f>���}�{�mA�G�+гn��dlb�
mX
�1�AP�|���(����qJ�%Ԣ�m�S'J��HZ"�M<���v?����;[L��+�iI� vз�>TtC�w��T���"�YA��wVg�]�W0�c�.]��w��$�:m��p� Ou������f�h�@�k���bһ���w4�*Q�"���,g��0Q����<� HUݜ���"��
����r��/�"�����^;j�yћR��u�p>���V����εXlxVHYEB    fa00     640�#9:���c�Ḿ�S�F��ђN����������֯+�������TdO�`�4gB��K��~�l�)p*�aS6�!�%s� '{�C�m�ڢ�g�x&�ٟ��1�m�T����TÔ�Cul��",h�+��T�wv������/G���}�%����hRҍkc��!�6A��o爉�F��c���חg��p�^�@��μ�gMɭd�9��G��ی�����e^T��Ŋ��2�()&1�M�t���s?���DÛ�Z�-TO�b��4���Ȯ�} [�gWRW^:44!a��c8�a���\a�XKX��I��7��W�������-�;�;ᢌ�Z�?��>����Kv�|h��� \�]���qs)����vg5�����)���A>�E�<_��._1û_pˍw�eAP�:/�Z�S�ۍ`�#{���c��^gZ=h�H�k�Ů*�rdX%�¿Ϛt���P�RSd;b��$�F�pt�"�\sG�>�-�1�ߖR�[;F^!����0F��yi��k��LǏ39g��k���I^7� �$.i>` ��Y��~�բ�-W�2��c��]s_��Z���o�?XR齭z��lJ�G̢�$V�^L!݂e?4�7μ�W��qF2�u����O&I�uZ���)���"����g7�H�`������¬����ʞw�8������"���ꗂU��oq�e5n������ �i�a��>�}�/����~KŒ�+]�V�s~/���%I�b�)�	�t�`;������u5��k_X��/� ��S��Qt"�|v��s�YV��}) ��%���e�V�
vR�p}�]X#f��d5A�B6
  �/��b	���-�PS��� �b��é}�T��\��'?�М�f��&aV�讝�_/1��"�BL�x*x�1{3b	�B�U[-��8�$!���5D�u�+!Ԁ�|� P�N_���re��!�]�u�NWjb3���9̓��&�1�W����<uf�m0�"]�� c��a�ƭO΋�=@7JD���>I׃lߟ���QgT�j�2?��#b���!ui5Ie��f�\�sy������;n���)�~��X���P�,(�
F�Q`�)ߓ�1(�2ٙ4�3o���<z@�@��n��
'm[׍ߺ��AƄa]�i���wTj/��Ǽ��c�Ey���|�a��+��Z��,}��>�z(�Z�n�p�tM�������9�k"ү�ӻ�����i�*=ޓ�:��L�ht�ߥفto�F��tS�2�����nJiM���s����C쏩;� n��,�b�dǞ�X��/[��s)��"��]���P���w���@��V��[l���~G�]�=�il��oM��r}!S�d/�o~�0U�:c��'��&����XlL*68�J�IF��dM�>�b���y��Wh���	�K��s�J����T�.vi^w��¾F&͸���,����9y��D-D?ؑ�r��o�c&�+�q��*��|����sH��e��'���C\"$1�y��V
����%ml��V��N�Oy'[=��sPW �KL�X����]R�3���"�rTXlxVHYEB    fa00     5c0�H0�.���,���P�Y>ER��҃� �`�����x+���ƴ��C 2���|��Q��u�}ł��.|^�'Pni;@u���xm;z��ݤ>�x�H�`#+'-PG�ir�.���qPã4�4s��7i)F�4m�^�4��G8;���~+C��j�Z���{��\n�q�A11����W��eiW��q�J��E?�wg�u�����"h�i=�۴<F˳�]o��7��
h���'p���ڊ�F��	��,��
	��K�k��j\V�FB��w�hBq�3Rx��"W5�5E��Cl��W߫�HŖ>�����|�S#� h���>�!�ז����e��RChXH��1�ܩ1�AZ��-�'���cyt�;L�Gl�>��GDw��yxku��6��J�2���B�a�r��0�_�c����[y�f�9w��Ӌ�,l:ҳuu�!I�]�OwXc��CK�!�ډ����y��hr�¼��&k�k�o��vu�sW�8	��C�Y�}���?d��S�ʣ e~*
�riV��rw�]���0g�ٿ-�#:��,���w�3>B��?�a����0�S{kku��M	Df�^���]���]Z��A�Jp^��c��v�,�x�C��+��=�� ��� ���/���ۺf6�B��+�?S�F% ��6�3��b�����~�*���� N1�����Z�ޗ����a/���>����ՁĘ'��t�����5�%��S8ok�v	p2h�����|�XS���ϊ4 ���,􇝀�_N���*~����
���ݞe����Z�XS�Bh����oú�{������:��B����T��<���&���aVbkh*����F:�$�$��6)	����r����x����C'~����J�������ev9`4ؕ-�,�c�G��$���f�C��J���@�j�o?6)ٽ1���|\�V=�ÒD)ǁ��w�Р�-��[����9��L/B�8I���U��QY��qg��܍̧�2)���<�aQH�^%�@�~�ZD]ni(�J�G��BWo��4��Եp�|��!��>D���WnX U(D7�ZA�����G?�D��q�d���׹n2��2��-��Ń�u�-�������}Q(���{���C�7�y���nx��Ķ�Y�ԍ�?�>>���w����<���+�����x�a+�i���_U��������̽ԁ���}��e�tDú@��_�%�^����'��^̌�Ob�==�&�ʉ#d{�M�nO'<� �t��_	m�n�pSZo�no���V��G&O�q9�ETt�} ��;;�G3w 5�Y���4ϕ��,R�)m��0����P��
RF'[k���C�Xe����E�3�� &��E��7��ĝV_�u��Ϧv2��Sߥm� �f]N}�����HX�\S�_lXlxVHYEB    d347     a90H�����݉��y�pw=˗��������m���5����i~��,����Q�H���� �]�	�Ỏ�E�z�@c�q�cM-��'���;y���C~������$�>,��b��� �Ҵ�.٘����������p��A���i��^�k�`jǺ_+��At�yR����,���+����Q����G�%�/���.�S�kO4���~��pd�E>{�����X�E�}�wB(ֈۆhZ����佨�n`'���	�U�~����Yjʋ�s��� �_~u��GnN���ȁe�H���?�#:�%<��y���NZ� �Ti݄g��!�FҾ�n�������L�j�w��A����\�"6D�C;#���I�+��S�F�[n�x��c�ۯ3�Ͽ֬-�w
�*D�Hoq���6E�`=N��`��չTG�`΅�`�:�˚��2�5|Pa�~�Փ_F$ͫ\1:�J�&��ẘ�f�>0!��r���~j�;I�x{WJd��u��O��O�5,�Hйmd7G,���#<��f
9�Z���[ϐ�/�S3��l� .'��*ꕟ`^eS�uȒ:�e����jB�L\y��y��ob�b��B~�\;�l��(�,4������T���dpD�uԵ�����1�t�R ��:��p�_1N<�`nk���H�u�Y�˷���wH5����??��ro_�S�m��D^�} ���i7;�*h0�1�rڈ�@.���#�Bk�q���KK ��,V���jI�t���������ng�(+�v���I�~���!嚯��Fz4��`�
D���ҩt�8����N�vϾ1Y*(�5j���E�����=8k����/�ߺ�Lr'�	�:�z�T<r�����S����b�q�՗̱��
�#빰�Z%~�r�Â�tX�+�����4�������m��v���Pg�𗏰�ݿ>�Oq
F��3|d*	&�'���K������k�Cm[��:j�B5_�S)_���>��Jī�H�.D���`�W��K�[��HgL��ۥ;Qy���?K ��@I]��/fud6�$\��Zꫮl���`Ҵ�����y����UB7�HQ����ƣ<pWnc�s䭸7@L��ݵ�OU~��R�.��ځF6���y����]d Ƀf.����AO"�v��Nڌ���ɃV6\��<�B����!��y��i,((��q�V;��(fSBVM��e}[���� ~� ���v]�^)�A
��K��2V���9��ߓ����V��^����M䈵�W�ju��'UCe�Y��Ѧ;���Ԇ�����_.��@��4�F�ף�l���W�c0U��dF���/)pG`���w�Φ�lC��*M�{뛉5*�z�bZ��x�텖��9W�����y �>:����R��AI�{<��+�iྋ�I�mG�aF#�)}��ؒ�2�3KɾÀ[Xr� ����O�-L��ϔS�O'T?t��\��yN
�M�Nj���5���%���a�^>r��'$�p���5�$��bF��~��)K�D�˒�K5h�s~�T��	RVT�y�Kwhn�\�4�@���;L/�Z�������06��Z, �.v�.�����<y���7~��#8��?�bST/�<�#�C�
+\�T!b=}����Γ�U��qz ����i���?Z `+���6�YI��qpu��ܕK�S����%0��դt������"��?huT�L�#l���P�@�1�'Xn+� [h���QQ��i-�N6����胅�ʆB#x�R���p����8�W��a~�|3q����e��_>��|rD���,0)}�5�S��m$]>؜|k� ��u�3�3�t�ׂ��<�����ȳ���'�`|����	�a|�C#�}ZQ�1��G+����z+�i"*���X)hx�n�`=�������t��`5�g@������s[|��vζ�B�/-��\�lέ�:�ǘ徂�ΘG�� ���t��=�`��M*,:�$�� rD� S0Ϙw(m���]���پ����ۆV������}o�O�@�&dd�~���}a-�sR�b��nn&մ�e �#��aRw�#���! ZcFj��c��r-�O�>h;$�ҧ�g��<%��:�]��F�6�F���㮧� ���	o8�-��y)�!>[�J6:f�ǁ� g*q�\�w��6Y�A�PJ�o"I>�_���O�~��Ϙ�{�kB#���ͺ���%&���1���vxQ^�i:�KO���1UU��&+�Ib�*�Z$s�V:M�DK���̫V��l92:��e�8�]��_z��ۊ�U?�����7��B��C��519��, $�廤��"��l,�9���[0��&;����^���e�g*c4��e���?/7Д�V��u�XC����n��rys��&��{ݪq�=}��y��ϲv��-R}�t���߉�)~�o�8*񪲝H���GYV�i�fQ��Adv_+��@VUGd��I�P`e���9Kq䨝�|�{uaG�\Wʷ	|0�Ο�����
�o�d��E)^�9�N��8yĶ���������&6���~�I�GX�����ںR`g7�"�o�u�
$������