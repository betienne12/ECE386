XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������+U1�[=�y3@����Y��U��/��$�1 �����`�d1Sr�k���Q�Ù�Q�kʃ���j��,{G��ih���d2��-������u��iS�\��^5����g��!��L�W�颡�ύ{�|������Y�� �>��,$�NcuA�\�U<����>u�wߔ)�"��m��Â���&Il��1c����U���*�j��sz��|��ϳvPP!�ɖ}Lҍ�޼�u��u4"
���bab��٢���3�Q�@�&_���v!'n�1�4m�����=go��6�#Ƀ�����阊�BBq&&���7��=�'���R���R����̱���Op��M}�(�4����j����lՍ]k�מ�@[@0Ӳ���토%���U���`e"ja�sK%�JtA����p�^*���V`ޏo��i!��y~U�!��.���u�:2�7a �dX ȳ�I��.���f�4V�E5����������O�{�qV�U\�������I6��1F�	*f
5�;���c~8�n5JuN�Bm�(��Q��wW�7�V�9fPyjl��x7�~��WO�IN�p�E��ZE�����ʁT���f��� ����ۮo�n��.ap��)E)���{�^��ɠ��?��iQʜ�3f���<ՃI����\|�t뤈M@�!�)�M>���������ʤ��;d�D��*��e�V���U�-o���L\��z���/� 0��ƫt6�;�8O�XlxVHYEB    1427     840�9[|wa�.Edϲ5�����ZġZ�������;l�\x��+4���1В�H�<;��l�xMyM����u��ה#���;ʚl~���¢y��S}�b��+{��Ou�X	�J�iqЁү\���?�����u��E��[��x+���:�F���É/7�'5�c�T��Y� ������c$�����{gZ�]��\���6���������q�'��oC���w2�i��Q^�����wh{�:��N���PoɊ����5a��~���Q�lĖ��uV�3RMg�2:��N�t�j֫���������j�`����8��u2�;��ʔ�{@�3P�\R�ۍ�>X�G��`��3)8L�[�����K��t���B�<CR&�ď!4�06ǎLK��r��9�8�떛N3���x}�FF$�Y��c#z�������
JP��z��'Ц^O%�.�ʍY�C�gO��X%��Fo���e�����e~.���Xs������4XYU�x ���c����,J�`$Ӭ��a��Q������{�x~L�s��߿a=�����Y2����f ,̈�U,���E�{k������ m%)(1Wm���?�N[�R(� ��~v@&����w��~x�LKܷ�j�!����@Nx��i?&.Ml�g����4�����D. n,��z��G�����@��]v���aL��Z0棷�Y���0���
q�f6���-�-���K���h�Ӡ���,#���Y�f��L(��hSv�6�zǸ���+�E:������Ji�u]�q����*��}d�<��Y�I�rK���p�/e����X�����BA��i7��[�4��&|��X��X��e��db؏x'�Q�����Y��o?��?��m>X*��s�by��^��nY��ۮ1x���0�#X�5��s;*���_g��Q�+�T��`m���I\w�YXD�$,P-��2����K���G6�-�K��t͏��*c8�|�vo�n>9�.�piLf��#v�8�Z�ws��a�X=o�b�!>A|���C��<�@
[pn.=b� ~����x|\L��,��0�k���4�(ӗ2>�BY�/�	�M�j#��c��+�.p}6'F*q!Q�CZB��_�g�*�j�ͻ�x�W_�X/ā�?5q��Qk�XJa�I��]��I�jc�X��q���¼���!�MNk��x����P;K�����[S��euXT��>�SwiC8�;�鞐^B��-Y^`���+�O��87����& �����@_�4���@���1B����%d�q���T����l��q�-�T=���w3�&g(;&�s\�n<��ik� �Cj�z����V<Ð��b)�^�k���Sҳ��~ ��#|�tiumO
�>�%�˚��+��y#�eA����p��TV%�|��G	��ң�u���j���(��6Y��:0�mr����N% {���ްу�uH���E+Ga�O��Ggr88y�}�!Rr�����chT�H/�qf��t��=�>@��be������{�ȳ~�_�<�����bd��x��8����\�O�CLOO?��K����³��<d��d�4�%���K��B�@�F�wlӠj����|�!^�wx �wCl(1[e���["���a�w�A ��/��6P��D{c̆�*�F%�ƹ��}@ƣڼ5�$R��ա Y*�V�o�Y6<�C��S���%��*�9��T��б��r��0r��9����`������8�V�0��mpw��+�$|h��*��(�� ����	}!��-2X[PMy��8O��Ӹ�Ϛ(�Nhp�����[�����X���UW��_b��+ >ͫ���fC-wu �:�i&�a�NM�\S)|��v<�&����~="�#�f�}��ɥ
|;+И��au�
f���bkR��F�(�s�Tԑ2���w��J���G����)��e��d�%enэ�el��R�=�niڙ�p1�F]0��������rm�t�E��\|@��9�����߻�����b��I�>tmY>"�$��l\�f��L�