XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_v�f ��NwT� 댏�MҰz���>����9�I8sS	�.�	ܛ�`UVF$_��9dI��u��Р�����|�wu��N�8^��9�Z�F����C�rH�͜�����t�-yO��P��#D�`��L·eu����D�߿e�C_��b��Qƿ%Q���a�P�Y�eH����a�;u�^��{�Zu��C �ܗa�Qg�<��RS�MZ�� ��\�+�$�m%C������y[�%;��N[-Y��������'��]��W�g���e�B��L2u܍3�trΰC�U��%x�.PH����h�r/��+1�n3PT�h�L�cN��������bY�JKړ�>�F�����Ⱥ��غC����fb�P�?�ҕ
�	+���^����{��pg!���g
*������ƬV{Q�A��<N[��^kp���Mb!��m�	��#a��D[!����ZC:�Q�69��,����E�G�ha��B~�Vul�̮P���ϭ~x��J� �QW��w�'V��������6G��j�6���8w�7�Ꮀ�
X�Ss�x �X"�T��"Y���OX'"�Y9S���j%��fMUǜɴO@�j���"5��ye��X�b�)���;a�cȟ�3<���1A	I<]����g��1j�$��iH���r���;��LA�.��ɭ�"�xˑYߑ`�Op�����c�%|E�Em�h�<������7N����2M�-W��G�T����?��6XlxVHYEB    fa00    2020Mo�*	���cvg�6�9B��t�E�L� e��U��h�~�7=���,(����e1��Z��Eu�)2��"��%ᇐ�Gt
�PbmC֏�CB�(���[�Gb��_ ����*��a��$����ܴ2D�� �D��w���E�ɜTy�#?
ʥL�!�R��?SWT���SFH���(����]�!�:�����C˾�W�����^!����>jӣ���t+@� ��c�XҬ\�����;�Lm�(g�qmֳd;mU��u�\�e��n�q��3�E��x�E����s_����l�Vi?7���X%;%h���/�֌:��K�59?+�E���l������?+1�dy���Pw`�y��i�����%���V0�j���7�r���F"_G�/��� n���PB2��x,�oԵQ�~�+��� ����!����,�E?Fp����.՟oa^7�S�.���kɕ�v,T��q���p���dx9��^��C�U:��P���9�S��t�KҎy��~,� rz�*�L�u��}����.
,Iz�`����Y�`o�33$�0	c���mv�����vy�G���rx��J��l
�E2!���f}�)�ևV�5�m��7B4�oi*rG����uU�
�,��rNzR�G4,*sѠ���oS!���]� a+G��k�Ĩ�'b�������@ĩ����Y�|َ�V	����W���q���wG�6� ���rV�x�������
��{
�mbS��z+�h{�;��2go�LJa�RK��G"눕�,�my@> ы,?����D�T�q��D��e��'�Usa��F�F�A�u�./�B�t;��c��MU)L:3�|�U.˼�!����$����z3֢�4Sx�Lk�6�L\�����
���I�|�,���>�p5�f�Ur}u�q����Gp�:�B�9�����x<��,S�9Y�a�|>j;�/D���i��>�Jv.c��l�����њ3�	�bEVms�}��X�/U�c� �jc�C-��<�� �!~|�v�SN��V�|x��cW�:��/ڏ)�*rz�����f��"p͋pe�A�0��5�m�W��,%Y0�qʕ"�2� ��Ha�М#_�Я������;��KoVCύ+L�43��`�����S���v���j�#F�k�F(v�D�Q���|�H(��:cA4��Z#��������;1DH��w��<Bk�2X�ȿ�Nb7<��zB%����I*I�۾��"�W����i��
c�;�mY�������*{:�,�pπ�ti�� ��s�1�kU��&�MU�D�夯�+,V�,1-n��$4YW{%`�O���Ʒ/�.�,I�xO[���l~��4�"�J���-#L��[�g���������	j�n��8q ����Q���9J��f�}`B4p�p �j�0��zĶ8�ljq�vS����q�(�9�6"i���Ph���ҏ�R�M�s���{��U�V��}(}�	x�$�A�g6�����:��b�{ *g�؂�kY��~��1y�Kj���\֝L��	ZO�lp ���*>ig�>J��/Jy��#�Z���S���;��\r[�gS:���5=:��p�J��^A��ÀnȺȦF[E��ĨK̕=�L%��d�1�i�ި�$��.�I �?P�C�,��;���ID��<f��/���ݗ۩�d�`|��^DXEj t8/��5���oDK�p�ɒ�%̵�mBj��2�ܩ� d-+�:����%JS�pB-H��F3�2 �4�VP���r�����(���z�O��@��e�eo��'<�g�?���x/�(O΀���nҊ;{{�pP�J�ɰ4���Ғ�Io}^$���KC��C�V����Q����S�dA�4ŉdI.C!��oӉ�k�Ӂ���{�X�VyG��@8�U���u�S���l�xq����*��26�m��&P]P}���Rx�tʎ�Tr����n�W�(n*;�#���R#?�im魹I{�U���ڷLc�ݙ��������Ԥ�n��J�0��.4r�.����Vr���I�>�W]�mK�#D�p,���qv��G���.$&TV`�&����S��w��k+s��3�i����(�\V��h6�m�pe�(W��3x��ә�2��$z^��d%�TȲD��9�:�Bb�=��[��K ���Dso�_O��m�C��6}t%�M���d��^/���ж�F�/����3��Y��f�wq�B�b�[잜�	���>� �j��q�w�2�k�tdd��KpMW�+�
f��$0�]��c��O)f�>�lV�#"R.k�u�zEw*�������	������k�|���k�X>ܕ91H�F^[k�-[�3���	۫����U�*sm�X�e~�"Zfi�u�I�����'��s���,�Wh�s=�w�]�`f�2�ٜ	�W�	v/~��{�ǥ&�qK���Xǟ*�:��
J|��A����%�7�vR����9��qj&����Q����!�Yd���<��:��wk2v|s��J�'�l5W��Gתw�u��ʬ��p���G�T<���M��l
��{��e>'/
+��\��n�1+g7U�O�@��ˆ�`������XR����jei���*�U-?QlƬV��������	��xT��f
ZkLN��0�$;3O �Z�����[��zB��A:*�����/�I R�����c�3^�w�Iӵ�Tsr�:��@f��|r�(�xz�Q���~��g����?�[����(0��Kd"ހ�ɛnؾ���(b�:��=�ZGc�}e���[
j����Ø�BL�0�MCWm��.���Ki���7��B8R慼R�fT),�K]鍿�$Y���~�������C|�%���<W���ye�{ԂHp�
�K*��A�9Jγa�-��I��2�0�h"��p�;!91Z 3GW�f&���V	���N�=�����X���kIj�Ts:��F�3ؑ��9�&:m���n4�u�<."�uXz[�U��	"�ױ#�E��<�_���.��`G�q���߹mf9IKL|��{'�jD]!�ȓRď���&�����T��S���jHQ�kh�e8�4�#�0Z�-�c�ER(�e��Q��|B�cB�1�9hRQ��<�F|i��S2���l���8"���@�+��|Tf%c�D��R���(��%�R>mL�6�������'�ϋ9�FF���n�$n�l]\�����"�%���$��6s��..9���'a��� DSV���OF��27N� _Cǩ�|�z�zz�搰�f�Ʋ�����pL�Z���I{>u�. �ם)A1�
6���QS�9�tj�X�3"�	�w��S��}凟�Uo�7��i�Y"x��4�y)�ޗ-°��5\�Sȭ��O�~����=2�5
	�uԬC�5OGPh;)H��V���<�	��%���7�쉖�Ś;	Y���G���D�ꃏ!ی��%�q�FR	�"�~+�����!`��WX����lz'����\�T�&���`?�r�Z����0Dž8 Z��S���m"�Б��Q��۾�Z��I%�y�L�Ž����ݳ�qn��P얢�����b���{�-��+�Śν}�w���,���� X������&1/�	\�^ӌ��Xz3�Z���7������IR�̊Ќ:�uY�E����j-�`�,{~�%�7chy�@MM�2���n�V�ֶ/�.B*}��df�K�+�^���J\��@�;��/4|���"{=�:����_ �j�}Fz�y�33�x#:�W'ǎH<m~J(��{�05#��mC�q��"��S������<)L�[c~��n����!�T��Ӷ��E��G�f�hƥz�ԚY�=�C��@�0�Ҋ]���7.��&Dx�p���r��B"ze��=��"��Z��6�M��;I�+�g�Ra]��ZՕ,��x�	V.��>O|^���A�sg>VnT�u�ֺ3�qv�4^e��^k��CMm��n��s��]о��r�d6�('�ˑ��X��̇���m�X�R\�{]��@U��F����3���ox9e�<�9\1晃�̢%��E4�f���d^U�IϪ쏅z��~s���!�6�-�)R\�QFԤ��� �*���0X��	za�9�W~L�r�0䳨C�=~��p��2��עa�Ω�|���M�P,Xá˹J'�	��Ӕ�^�������Z8�G�vA0�c<����L���8X��ưc^��m�dГ�t1c���@��[��y�)";2Iz�bv���=��M������$&�&����+,q(3Eo���.�YKu��G9Yk!8׌j��A �~���RS��<��d�JU3���%��� @2`�f$�B�5��o]���-���ώ�:�J�UM}�������w�6�~ht�~Yq��:t�^�p
/�7������E�1�Kv)��E*��s"�������Q�bc�4�����%�%_�0n"~C˾=[Ԉ3\ٍ^nߗ�� 1�r�����Œm^��� CЩH��������_���]cc�f�� M�~�~���@�rK̷�17������BH\�����V�xpM�lF���=H��P����I�L����0�{]]��9���ٻ��Ȃ<��!C�E��G�������}��P 9�����Y<�wh����)��D���=��R�|�� ��\����B�+q��:���Z��Ĳ�����/���p���ۦ�3� aBb6d.#j�ܔ��F����2�I��<?�rœk�$�a�U9L>9�.���h5x֟�3����sT"] ��(��o��B��0S��?�}Ͱ?��k�2��	sv������-f0���N�]�8���T�W�ŭ䪝^�<I=�i������~�W�i��1JdK�k�2(g�P�Y�r�ܽw�S,:�E��/a7q���
�L:gBn|�G�*���u��.��]�&5�k8h!3H��1�-x��v=��pd`��#�l���#]��즊��T�8�~š�A~�O�=���)F\�P�{(����5������X��/��h�� ��{wbXc�l*��y���&]N��H#���K,�z	<{�+7�/��	�
�vj5Brf�k1�X���(F���h�����R�M?�8�wN$)>nTp����U���̼�,	��tr������������	����짙B�iE�| ��l���v3X\�B�u�\������S�Pg)X.����Y ���WG�A:�I��CNr�Л���͵x��GH<�JaQ�lȿ�$R!s��'d���e�� ���⇞u�IU��1�}K�}�ͩ�(�F�U��^�����
Sm��ۼ*�-�ؘ��ra�e���&�~BL�K���
i��F�vh��?�z^
$CF�Sy�e�]��� ��@�"D?b$��#���P3�R[&��tLy����u����g���&���_<�.K�'@�/�`u`-�@X�3��6�1���T��.&���v]:�V�����,�)���:����P�r�zHB��[�����\�ŕ�Y�
/-��[Qkz�V$�֧�$���t�el�"R���$Й <�������H�1�U8��vg��J$�|�`�Z����.�3��~r�'/�R��,���0�8�4=�����?�C��G����E����%x����T��X� �`D��lG�g=������E[�"�������v�O��Pi`[��(��ƴ��V�r�i�7�r<�W,zr��B.�M������#�4J�N[��,�8�+�xYzhn%����xax�^hCgy�	X� v�W�[�#�8QXǜd�fu�O�*(�xS^�3����V����� ��8V��:t=�;gd�D>��ù����d�R��E=#1Ry�[�_wQ�L�y&���̓���iڥXD��ʢ2��72<��k%�; ��;��

Ή���Nk��wP�s�ہ���D?�B�6A��`�Wbk�-G"�+��@c���w� s��T;cJ�!��������q,P��˯��n�t������(�@�)EA�tR����F�`nl"���)�9Xx�(�w8�ϝ���}pV�|\�qZb���3brd��+2V��E�M�{����E�`M��)���FS0_�#�"��A�;�*�b�ӟ�cJ:=|̝`ᮻn�*\O"��yM���	�U��:(&|��W|���/�f*��(@�5��b���%�F�BT���	���֥�����f�7`K�(�x��p��N�tm�i���1� �u�n�L������ˆ� ��C�E~)3��u}��Zh�у��� ������\����dIvKD�^N�X3�����Z�sP�߇�}��P���{i���uj��I�^I��?�|*RM+�]��@��zh�#jPA���X�ܽ�0�	��FF�1�v�)����>Y?*��j�m��'-�mYHiO���> ЈD�K��*N!k�!m�!�
��pK`O�ew7�v0&ƾ�gQ�c g�<��L�HsF�Fv�aL�Zp�H���/��A�\�N�,yx�(���|..�t���y����Ի�Lܟ�	x"�ၘ��c$�?�^x����'//|���ͫ݀���+�m-Th;����6Lf�}�
=�o���Vm�D��2h��
)FiG���s�)M(���G!�C�'>c�5��q�)��� B�s��BgVB��_g
q��L��׎񠥚݃�C�q�>WTp��q� �M��ٖ�����v�����vNьd�v��*�?Vk
%�����m�$�'H�"7�R�ĺOcZǩ柤v���J��dȘ�U[��fa"���#?�#I(��{�8ݏ�9�6�.y���X1e�a���W*�u��D^<]�HZ�ڠ�g����q}��2?�ވ�Jz�$R
?Q��-�fA��i�*|��,%i�LP�U�%��o<���Wdr�8mK+�4��*b��ƣ;���-��	�43�����\Vo�2�=5��)�zKo�
RM����%�t�<(�Av�
�A&rur�IS��-N�۠A��X�;7\����2��o�Z�������]K^5�Eo�
���cFB��d���P{D=�p]��	u�R��k7��	��)B�m�Zw/�G^��~�6d%�����K>Ir\��+�a}C$_���[��4��mAҙ������ZXw@_�Sx���k�����,�47L�vy�����;p(�Zŀݿt����m\���<�O�} 4�d Q�"j}cW�)��Ő}$�;A��enlb�auF�(BC�d�g!)���0pr�X�����l�h�IE��*�I�S�ޙ!�A`���nC�O=���zQm7J�WȽ�&��5&�e1b�%��Ǩj����zM��{�׏�/�ސv�I�Fj�O�;���W���h������������7�]�؅qnR`6ý#�= ���3�w�hR'H�g��	̈́n+X��JN�yk��6$�j:���Y�u�e������` #'1���z�m��sl��h�������3yֱaB�M}����d<���tB�V�Ÿ�$,j1:y!���w�e�XT�-��G��04L3�c^>��z���Kl��a�J��'�n�x����-����eP�!P��?"U��Va�(i�{K���fe�)Ֆ��B[��W��$L8%R-�1�E�6i����q�z�)r(x��D��GAi�Ǿ�k��Vm�.���p�8��x^S%�d;��3:�Yw���cNt�v9
�SS� T�T�����ȥ�����5ݠy��=}U͕ B,�r%}�ߊϠ�Oo�Htn"]R�Ӽ��ƕKۣo��gy��R�U�]x����=J-�Y_ˢ��$���ٲ��)��
��V@��>N]���j.i�����x�O�*t)nۀ����+LI[g8��g%<hK �HTÕՓ��F*�Pt͏�>�쨺��7�u�}b%�v������[~����&]+!�Vf#XlxVHYEB    cb82    12b0�wL���W�	�~'ɣa<e�/5<W�	��c?��Pr�{z�J��������6�I�ːó��[L$��K��vi�![��6���R�u#�x$ݾ�b�l����M)����L�²���I��K�k�]@޽_I��d�Ez��(x��W�y�{ ��,r5J�X���"Khşo��8$C�3W ����S�ҷ�9hF���F��W���g��c���3/�7qݬ��ͬ����*���ps��X#L��h�Py���"C�'A�%��؏��+���m�Szc��9G�T�,_N��D�V�_��u������H�t/�;O]t:�V�L1t�7 � U@�¢�)�ǀ	O�'��ȯ��u*�R���e9�`\2�G��N��+�",q� �w({����
cʎu�`�L ��YBvM+�큶�k�fڇ�Ձ��_c4"���U]���h���s��N��9^��Ap.�����Y%�ÿ2_��;5iXG��5�
M��e(�m�f�_�"O��ғ%�uO���y��k�>������U{=�}�IBpR�K���[P��<�r�f�#���� �=�va��*[~���G���1�ZJa�3%z��x��fk�1��V����E�r�V�*e[ˡ�S]��X��DoM��|����`�������_xJi�GR�/��waǢ%��G�5��2I�A��E]��k�V�t�_O��\Y��y����ЮD�u̙�i�o Hk�'��fV�� ��*R��1���uC[o,<
_;Ţ��!rz�������FjC��ߎ�9v����'�\��(�o#��)i؛ �\t����Zp/��!+YwnIm��̈́e"D�nU\�`�3��y���R���\�uS���~`���ZP��|�>7�x�6p��ʙ.@��D3��!�U�8�)iN^ڤ�T)7�F+q�wDi�UD��P��>dJ���n�2�����y�������&���#0�7�bfSc֌��1�)��mK���}��ޗ��?ݫRZ8_s��B V���Ҵ�Q9|R[u7����KwH 1#��8���d����PN�\t�Ӥ��OC+��罶f�r\Q��_�dv�-rg�ݤun�6���dp�u�G���_JY��qS���9��HJ��U��fqm�Ʒ3� b������+@`��~�?�;�x�
&��_��R��PObb�n(�O�����y�Kb�_u�v%�)$�գ�(�@ȇ��Dz�TE=]QΤ���h����^�� ����VxWʖ��u����e3�·g~�r([����*q�Gwf��f\6�<@ x�x��n_ٰ��]�1�H�YxJ'�[ �:�h��/�[�@�ۓ*Q�]���IG�AGV�7,�����e��[aR�[hۯ�&�9��"��><e�6.u�
+�I�Bެ �^�JT����B0:��nU�fg��0#,2-� _̵�p�� ����GEE5*�5���;�8}�8(Ϫ*T��A�<ɦ!���4�������12hM����c�6:H����@�w*�&��e@ �������?	1�Xē\���5-B��%d�4�-H%f��Ԇ���H���r^+}Ȓ`XX�n�cS��A ot�d0U�b�p�/m��� X�,F\�:�+/
IM����3�|�[��7��,�Q���*s~��(|}��Q����0�M�`q -�S�s9��$5����7X?;�o��1���9��^��1��q�c/.��Ru1��0�92}C�e���_i���%�<!+p�L+|O7Sn���o�j�JZ��鱭��ʿ���Y;<��H����A�~�kn�ޝ��*ڼg.wN�[�U�"nJ�/:^�*��2���4V����L��E�)�&��!z: ���|L���8��|�k���I"}��+�0�-�W|���d�����w��	"U7���@���!p�VeLE�%� �5kI�M����o�/27��cN�3cYa���}��-�$T��@�ᘭ5��3pi�T�xx��ף5����� ����^��_24�[�.��o�_@,lDP���~�,��9�ŹV��J�w�4����3Ů(��]���?y��Z.$�d�W���E��pj��������꯽�I[��kYrd���ě~��t� ���G��ߥ$gW�����$Z��z��7�'�78�\�\]���򢓑LDr\���W޶�����c��8��c�=�K}�K�{�n`�����Í����� ���=̰�E_:Ѳi���V�R d!,�¨!�!�0�[��`�!T�.�z���$�-$��w!y}��ȣ�������L	X�wg�0V�((�z2�:�zH�s'�;G��7�"�9�J_���ᷯw��Y�-�ZLU3îGt�[M��#����lT����ӛ�L�Z.�$e+�]W�����Xn�2�X�qܻ�n�o0�w�0X��Y���N��f�Q��n����m��>!Vc5˪P4;f��W���`�X\m! o2�o}Ѩ�?l+:؅��C$��\��N��غ.�&k����7j�Ia uՍ+������Q����ǅ�I�j!�8g�_/�>F�3qH��/����� ����
%dQak�Zz�Vb��_e��~q��7fii���<�{�� �$�Q�e�i��@�;H4�	���1�Q ϗU�ؐ"榌�"�7TR�~����)W��a*�I�5u��S�'e�?`v#��@ۍ<ɟ"-v<ݪ���-���J�f��v6`"�S��j.�P����M2|6�����,���B���m�s�����3�qf1��T�d�Eag�U����L�|9��=��dJ���:�D�0Z�"8���y9=~I"�x$}h�e�=�_Ɯ�+-�^2}5�g�.�oH����ge>9���a��z#���h`畔Gt��k�l�V̛|�ǵ��2�4�����}N�b?
�up��7�p�*A��h���A$")��#�g�������k|����D2j?zC
�+ۏ[��4ڑ�f�B��O*���,��u�̙�˜���^>��lS���}���9o�6J��=X$�l�.��X���g8��M�Q'���ت:�0�y��p)ZV��|7��V�M9mͥ�ܗ_���
�=��bk��v��Sۛ�Z^��Ek���I�Ƈ�с��I���X>)�1��&�7�L��s\H�8{���3 �G���:N�>֪����(c{d�'��]��y~8���\�O[�[�ֹ_�50�n	���w��0�z�Aq{jG.�M�L=
 ƚ�Z�`��ޟy�L^�<y(�kz��2��HT�r$�?"��"�ϛ�K�_4(���dz5��MTξy eVYh B�>I�M�e�2=�M�EX~3��J��ٶD#
�'�x,Wi��W�!	�$�=�4E��:�m���W�����pn{��ZaΓ�:�p��W)b�<�*f ��}w�t����Ǟ��}�O�t6�'L�ec�@�K��E���=���G�y;"�m/�F���eV��A�m�/�n�z�J��?��L�0�<'�"^���շ�Fݾ����� �)#$iIt�/�})|���	2�E5#�إ��}~�8�ٙb>8ტ��S��>y�,4�x(�ƫ;Ǖ
w��y{�;�+���=��n�dnA�zsc����w�d��4G����D���F>��(İЎf�.d���'�z�[�Ѡ���9u�$���~:
���^M����ϵe��?YruzW&���R8̼>�ze�$�NK�~���Ip!���"1�(ؒ��	�m�-!	��W�E��4�Mxcs ���@�	��g<�%� ڔ�g���uAN )dIͺ�y�ъm��7����U��j�S����_K��Q����2���wDx���.�K����gX���:����ȏ��ݧ��g��]�J�˂���2�Ͱ�����w0��3;�D�a��stB��m-��9�i=��aR�E��GӶ}M���	6�4L�|Y��6~�/>�.Y=�RC+�Pb��-J�����&��9����~�*j{�bضҁpK�/�?'!ogbu(��I[�ΰl�}��	3gJ\�2pU����4������6��#�S��9� t����x�y�ҒQ��C�-\ѴZR�r|\y������PIb�l|�Dq�bc���[/
���-�Ȭ�D�TK;�����,8�Y�5��>�i�K!�}�Y��f�g�ݫB�K/�o״�~�.R���ݔ+���'�cԇ�����Z,'!Ga�a������͏U6e_Y}~\� zjI��BJw�Lf݌�Wz/��g���_p����Q�[�!j�F��1�7N�1ً���� �A�9���:S�$�;p��́�c� �������)�� ( �����+��� �ȽX���L�	�@TH`�?�*�/���D�H�gf��	)X${�pNW��v٘y����Kl�������k��^<7bl��{Ә��%X6|�˸��ў�os]���i�ʾɘ�̵����A�-��4��`�4�@v[����{[�Ϲs͟>��ʹ0	%s�3���_:�"4����q��M\�ty/h
�����	��s�K��rϙ'��7���s���¦����~N�=�M� r��ݱ��YXC�`���5�JE3\2��R�w��~�焹ҪOXH2w�AR���B���<8֛��f,��`W	�p��*|�